module FullAdder(
  input   io_a, // @[src/main/scala/dadda_tree_mult.scala 6:14]
  input   io_b, // @[src/main/scala/dadda_tree_mult.scala 6:14]
  input   io_cin, // @[src/main/scala/dadda_tree_mult.scala 6:14]
  output  io_sum, // @[src/main/scala/dadda_tree_mult.scala 6:14]
  output  io_cout // @[src/main/scala/dadda_tree_mult.scala 6:14]
);
  assign io_sum = io_a ^ io_b ^ io_cin; // @[src/main/scala/dadda_tree_mult.scala 14:25]
  assign io_cout = io_a & io_b | io_b & io_cin | io_a & io_cin; // @[src/main/scala/dadda_tree_mult.scala 15:46]
endmodule
module RippleCarryAdder(
  input  [62:0] io_a, // @[src/main/scala/dadda_tree_mult.scala 32:14]
  input  [62:0] io_b, // @[src/main/scala/dadda_tree_mult.scala 32:14]
  output [62:0] io_sum, // @[src/main/scala/dadda_tree_mult.scala 32:14]
  output        io_cout // @[src/main/scala/dadda_tree_mult.scala 32:14]
);
  wire  fa_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_1_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_1_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_1_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_1_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_1_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_2_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_2_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_2_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_2_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_2_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_3_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_3_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_3_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_3_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_3_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_4_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_4_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_4_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_4_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_4_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_5_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_5_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_5_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_5_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_5_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_6_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_6_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_6_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_6_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_6_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_7_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_7_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_7_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_7_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_7_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_8_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_8_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_8_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_8_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_8_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_9_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_9_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_9_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_9_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_9_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_10_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_10_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_10_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_10_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_10_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_11_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_11_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_11_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_11_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_11_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_12_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_12_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_12_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_12_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_12_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_13_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_13_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_13_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_13_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_13_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_14_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_14_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_14_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_14_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_14_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_15_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_15_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_15_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_15_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_15_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_16_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_16_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_16_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_16_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_16_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_17_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_17_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_17_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_17_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_17_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_18_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_18_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_18_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_18_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_18_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_19_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_19_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_19_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_19_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_19_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_20_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_20_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_20_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_20_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_20_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_21_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_21_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_21_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_21_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_21_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_22_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_22_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_22_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_22_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_22_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_23_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_23_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_23_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_23_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_23_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_24_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_24_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_24_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_24_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_24_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_25_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_25_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_25_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_25_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_25_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_26_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_26_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_26_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_26_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_26_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_27_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_27_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_27_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_27_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_27_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_28_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_28_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_28_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_28_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_28_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_29_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_29_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_29_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_29_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_29_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_30_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_30_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_30_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_30_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_30_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_31_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_31_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_31_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_31_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_31_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_32_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_32_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_32_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_32_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_32_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_33_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_33_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_33_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_33_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_33_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_34_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_34_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_34_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_34_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_34_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_35_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_35_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_35_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_35_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_35_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_36_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_36_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_36_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_36_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_36_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_37_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_37_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_37_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_37_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_37_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_38_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_38_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_38_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_38_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_38_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_39_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_39_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_39_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_39_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_39_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_40_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_40_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_40_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_40_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_40_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_41_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_41_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_41_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_41_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_41_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_42_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_42_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_42_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_42_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_42_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_43_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_43_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_43_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_43_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_43_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_44_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_44_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_44_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_44_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_44_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_45_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_45_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_45_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_45_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_45_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_46_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_46_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_46_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_46_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_46_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_47_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_47_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_47_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_47_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_47_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_48_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_48_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_48_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_48_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_48_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_49_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_49_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_49_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_49_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_49_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_50_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_50_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_50_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_50_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_50_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_51_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_51_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_51_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_51_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_51_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_52_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_52_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_52_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_52_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_52_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_53_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_53_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_53_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_53_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_53_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_54_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_54_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_54_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_54_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_54_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_55_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_55_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_55_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_55_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_55_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_56_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_56_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_56_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_56_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_56_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_57_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_57_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_57_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_57_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_57_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_58_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_58_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_58_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_58_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_58_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_59_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_59_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_59_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_59_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_59_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_60_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_60_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_60_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_60_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_60_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_61_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_61_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_61_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_61_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_61_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_62_io_a; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_62_io_b; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_62_io_cin; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_62_io_sum; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  fa_62_io_cout; // @[src/main/scala/dadda_tree_mult.scala 49:20]
  wire  sumBits_2 = fa_2_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_1 = fa_1_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_0 = fa_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_4 = fa_4_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_3 = fa_3_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_6 = fa_6_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_5 = fa_5_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire [6:0] io_sum_lo_lo_lo = {sumBits_6,sumBits_5,sumBits_4,sumBits_3,sumBits_2,sumBits_1,sumBits_0}; // @[src/main/scala/dadda_tree_mult.scala 59:21]
  wire  sumBits_8 = fa_8_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_7 = fa_7_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_10 = fa_10_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_9 = fa_9_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_12 = fa_12_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_11 = fa_11_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_14 = fa_14_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_13 = fa_13_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire [14:0] io_sum_lo_lo = {sumBits_14,sumBits_13,sumBits_12,sumBits_11,sumBits_10,sumBits_9,sumBits_8,sumBits_7,
    io_sum_lo_lo_lo}; // @[src/main/scala/dadda_tree_mult.scala 59:21]
  wire  sumBits_16 = fa_16_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_15 = fa_15_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_18 = fa_18_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_17 = fa_17_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_20 = fa_20_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_19 = fa_19_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_22 = fa_22_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_21 = fa_21_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire [7:0] io_sum_lo_hi_lo = {sumBits_22,sumBits_21,sumBits_20,sumBits_19,sumBits_18,sumBits_17,sumBits_16,sumBits_15}
    ; // @[src/main/scala/dadda_tree_mult.scala 59:21]
  wire  sumBits_24 = fa_24_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_23 = fa_23_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_26 = fa_26_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_25 = fa_25_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_28 = fa_28_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_27 = fa_27_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_30 = fa_30_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_29 = fa_29_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire [30:0] io_sum_lo = {sumBits_30,sumBits_29,sumBits_28,sumBits_27,sumBits_26,sumBits_25,sumBits_24,sumBits_23,
    io_sum_lo_hi_lo,io_sum_lo_lo}; // @[src/main/scala/dadda_tree_mult.scala 59:21]
  wire  sumBits_32 = fa_32_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_31 = fa_31_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_34 = fa_34_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_33 = fa_33_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_36 = fa_36_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_35 = fa_35_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_38 = fa_38_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_37 = fa_37_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire [7:0] io_sum_hi_lo_lo = {sumBits_38,sumBits_37,sumBits_36,sumBits_35,sumBits_34,sumBits_33,sumBits_32,sumBits_31}
    ; // @[src/main/scala/dadda_tree_mult.scala 59:21]
  wire  sumBits_40 = fa_40_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_39 = fa_39_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_42 = fa_42_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_41 = fa_41_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_44 = fa_44_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_43 = fa_43_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_46 = fa_46_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_45 = fa_45_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire [15:0] io_sum_hi_lo = {sumBits_46,sumBits_45,sumBits_44,sumBits_43,sumBits_42,sumBits_41,sumBits_40,sumBits_39,
    io_sum_hi_lo_lo}; // @[src/main/scala/dadda_tree_mult.scala 59:21]
  wire  sumBits_48 = fa_48_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_47 = fa_47_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_50 = fa_50_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_49 = fa_49_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_52 = fa_52_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_51 = fa_51_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_54 = fa_54_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_53 = fa_53_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire [7:0] io_sum_hi_hi_lo = {sumBits_54,sumBits_53,sumBits_52,sumBits_51,sumBits_50,sumBits_49,sumBits_48,sumBits_47}
    ; // @[src/main/scala/dadda_tree_mult.scala 59:21]
  wire  sumBits_56 = fa_56_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_55 = fa_55_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_58 = fa_58_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_57 = fa_57_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_60 = fa_60_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_59 = fa_59_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_62 = fa_62_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire  sumBits_61 = fa_61_io_sum; // @[src/main/scala/dadda_tree_mult.scala 45:21 54:16]
  wire [31:0] io_sum_hi = {sumBits_62,sumBits_61,sumBits_60,sumBits_59,sumBits_58,sumBits_57,sumBits_56,sumBits_55,
    io_sum_hi_hi_lo,io_sum_hi_lo}; // @[src/main/scala/dadda_tree_mult.scala 59:21]
  FullAdder fa ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_io_a),
    .io_b(fa_io_b),
    .io_cin(fa_io_cin),
    .io_sum(fa_io_sum),
    .io_cout(fa_io_cout)
  );
  FullAdder fa_1 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_1_io_a),
    .io_b(fa_1_io_b),
    .io_cin(fa_1_io_cin),
    .io_sum(fa_1_io_sum),
    .io_cout(fa_1_io_cout)
  );
  FullAdder fa_2 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_2_io_a),
    .io_b(fa_2_io_b),
    .io_cin(fa_2_io_cin),
    .io_sum(fa_2_io_sum),
    .io_cout(fa_2_io_cout)
  );
  FullAdder fa_3 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_3_io_a),
    .io_b(fa_3_io_b),
    .io_cin(fa_3_io_cin),
    .io_sum(fa_3_io_sum),
    .io_cout(fa_3_io_cout)
  );
  FullAdder fa_4 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_4_io_a),
    .io_b(fa_4_io_b),
    .io_cin(fa_4_io_cin),
    .io_sum(fa_4_io_sum),
    .io_cout(fa_4_io_cout)
  );
  FullAdder fa_5 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_5_io_a),
    .io_b(fa_5_io_b),
    .io_cin(fa_5_io_cin),
    .io_sum(fa_5_io_sum),
    .io_cout(fa_5_io_cout)
  );
  FullAdder fa_6 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_6_io_a),
    .io_b(fa_6_io_b),
    .io_cin(fa_6_io_cin),
    .io_sum(fa_6_io_sum),
    .io_cout(fa_6_io_cout)
  );
  FullAdder fa_7 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_7_io_a),
    .io_b(fa_7_io_b),
    .io_cin(fa_7_io_cin),
    .io_sum(fa_7_io_sum),
    .io_cout(fa_7_io_cout)
  );
  FullAdder fa_8 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_8_io_a),
    .io_b(fa_8_io_b),
    .io_cin(fa_8_io_cin),
    .io_sum(fa_8_io_sum),
    .io_cout(fa_8_io_cout)
  );
  FullAdder fa_9 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_9_io_a),
    .io_b(fa_9_io_b),
    .io_cin(fa_9_io_cin),
    .io_sum(fa_9_io_sum),
    .io_cout(fa_9_io_cout)
  );
  FullAdder fa_10 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_10_io_a),
    .io_b(fa_10_io_b),
    .io_cin(fa_10_io_cin),
    .io_sum(fa_10_io_sum),
    .io_cout(fa_10_io_cout)
  );
  FullAdder fa_11 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_11_io_a),
    .io_b(fa_11_io_b),
    .io_cin(fa_11_io_cin),
    .io_sum(fa_11_io_sum),
    .io_cout(fa_11_io_cout)
  );
  FullAdder fa_12 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_12_io_a),
    .io_b(fa_12_io_b),
    .io_cin(fa_12_io_cin),
    .io_sum(fa_12_io_sum),
    .io_cout(fa_12_io_cout)
  );
  FullAdder fa_13 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_13_io_a),
    .io_b(fa_13_io_b),
    .io_cin(fa_13_io_cin),
    .io_sum(fa_13_io_sum),
    .io_cout(fa_13_io_cout)
  );
  FullAdder fa_14 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_14_io_a),
    .io_b(fa_14_io_b),
    .io_cin(fa_14_io_cin),
    .io_sum(fa_14_io_sum),
    .io_cout(fa_14_io_cout)
  );
  FullAdder fa_15 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_15_io_a),
    .io_b(fa_15_io_b),
    .io_cin(fa_15_io_cin),
    .io_sum(fa_15_io_sum),
    .io_cout(fa_15_io_cout)
  );
  FullAdder fa_16 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_16_io_a),
    .io_b(fa_16_io_b),
    .io_cin(fa_16_io_cin),
    .io_sum(fa_16_io_sum),
    .io_cout(fa_16_io_cout)
  );
  FullAdder fa_17 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_17_io_a),
    .io_b(fa_17_io_b),
    .io_cin(fa_17_io_cin),
    .io_sum(fa_17_io_sum),
    .io_cout(fa_17_io_cout)
  );
  FullAdder fa_18 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_18_io_a),
    .io_b(fa_18_io_b),
    .io_cin(fa_18_io_cin),
    .io_sum(fa_18_io_sum),
    .io_cout(fa_18_io_cout)
  );
  FullAdder fa_19 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_19_io_a),
    .io_b(fa_19_io_b),
    .io_cin(fa_19_io_cin),
    .io_sum(fa_19_io_sum),
    .io_cout(fa_19_io_cout)
  );
  FullAdder fa_20 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_20_io_a),
    .io_b(fa_20_io_b),
    .io_cin(fa_20_io_cin),
    .io_sum(fa_20_io_sum),
    .io_cout(fa_20_io_cout)
  );
  FullAdder fa_21 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_21_io_a),
    .io_b(fa_21_io_b),
    .io_cin(fa_21_io_cin),
    .io_sum(fa_21_io_sum),
    .io_cout(fa_21_io_cout)
  );
  FullAdder fa_22 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_22_io_a),
    .io_b(fa_22_io_b),
    .io_cin(fa_22_io_cin),
    .io_sum(fa_22_io_sum),
    .io_cout(fa_22_io_cout)
  );
  FullAdder fa_23 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_23_io_a),
    .io_b(fa_23_io_b),
    .io_cin(fa_23_io_cin),
    .io_sum(fa_23_io_sum),
    .io_cout(fa_23_io_cout)
  );
  FullAdder fa_24 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_24_io_a),
    .io_b(fa_24_io_b),
    .io_cin(fa_24_io_cin),
    .io_sum(fa_24_io_sum),
    .io_cout(fa_24_io_cout)
  );
  FullAdder fa_25 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_25_io_a),
    .io_b(fa_25_io_b),
    .io_cin(fa_25_io_cin),
    .io_sum(fa_25_io_sum),
    .io_cout(fa_25_io_cout)
  );
  FullAdder fa_26 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_26_io_a),
    .io_b(fa_26_io_b),
    .io_cin(fa_26_io_cin),
    .io_sum(fa_26_io_sum),
    .io_cout(fa_26_io_cout)
  );
  FullAdder fa_27 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_27_io_a),
    .io_b(fa_27_io_b),
    .io_cin(fa_27_io_cin),
    .io_sum(fa_27_io_sum),
    .io_cout(fa_27_io_cout)
  );
  FullAdder fa_28 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_28_io_a),
    .io_b(fa_28_io_b),
    .io_cin(fa_28_io_cin),
    .io_sum(fa_28_io_sum),
    .io_cout(fa_28_io_cout)
  );
  FullAdder fa_29 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_29_io_a),
    .io_b(fa_29_io_b),
    .io_cin(fa_29_io_cin),
    .io_sum(fa_29_io_sum),
    .io_cout(fa_29_io_cout)
  );
  FullAdder fa_30 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_30_io_a),
    .io_b(fa_30_io_b),
    .io_cin(fa_30_io_cin),
    .io_sum(fa_30_io_sum),
    .io_cout(fa_30_io_cout)
  );
  FullAdder fa_31 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_31_io_a),
    .io_b(fa_31_io_b),
    .io_cin(fa_31_io_cin),
    .io_sum(fa_31_io_sum),
    .io_cout(fa_31_io_cout)
  );
  FullAdder fa_32 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_32_io_a),
    .io_b(fa_32_io_b),
    .io_cin(fa_32_io_cin),
    .io_sum(fa_32_io_sum),
    .io_cout(fa_32_io_cout)
  );
  FullAdder fa_33 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_33_io_a),
    .io_b(fa_33_io_b),
    .io_cin(fa_33_io_cin),
    .io_sum(fa_33_io_sum),
    .io_cout(fa_33_io_cout)
  );
  FullAdder fa_34 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_34_io_a),
    .io_b(fa_34_io_b),
    .io_cin(fa_34_io_cin),
    .io_sum(fa_34_io_sum),
    .io_cout(fa_34_io_cout)
  );
  FullAdder fa_35 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_35_io_a),
    .io_b(fa_35_io_b),
    .io_cin(fa_35_io_cin),
    .io_sum(fa_35_io_sum),
    .io_cout(fa_35_io_cout)
  );
  FullAdder fa_36 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_36_io_a),
    .io_b(fa_36_io_b),
    .io_cin(fa_36_io_cin),
    .io_sum(fa_36_io_sum),
    .io_cout(fa_36_io_cout)
  );
  FullAdder fa_37 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_37_io_a),
    .io_b(fa_37_io_b),
    .io_cin(fa_37_io_cin),
    .io_sum(fa_37_io_sum),
    .io_cout(fa_37_io_cout)
  );
  FullAdder fa_38 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_38_io_a),
    .io_b(fa_38_io_b),
    .io_cin(fa_38_io_cin),
    .io_sum(fa_38_io_sum),
    .io_cout(fa_38_io_cout)
  );
  FullAdder fa_39 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_39_io_a),
    .io_b(fa_39_io_b),
    .io_cin(fa_39_io_cin),
    .io_sum(fa_39_io_sum),
    .io_cout(fa_39_io_cout)
  );
  FullAdder fa_40 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_40_io_a),
    .io_b(fa_40_io_b),
    .io_cin(fa_40_io_cin),
    .io_sum(fa_40_io_sum),
    .io_cout(fa_40_io_cout)
  );
  FullAdder fa_41 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_41_io_a),
    .io_b(fa_41_io_b),
    .io_cin(fa_41_io_cin),
    .io_sum(fa_41_io_sum),
    .io_cout(fa_41_io_cout)
  );
  FullAdder fa_42 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_42_io_a),
    .io_b(fa_42_io_b),
    .io_cin(fa_42_io_cin),
    .io_sum(fa_42_io_sum),
    .io_cout(fa_42_io_cout)
  );
  FullAdder fa_43 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_43_io_a),
    .io_b(fa_43_io_b),
    .io_cin(fa_43_io_cin),
    .io_sum(fa_43_io_sum),
    .io_cout(fa_43_io_cout)
  );
  FullAdder fa_44 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_44_io_a),
    .io_b(fa_44_io_b),
    .io_cin(fa_44_io_cin),
    .io_sum(fa_44_io_sum),
    .io_cout(fa_44_io_cout)
  );
  FullAdder fa_45 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_45_io_a),
    .io_b(fa_45_io_b),
    .io_cin(fa_45_io_cin),
    .io_sum(fa_45_io_sum),
    .io_cout(fa_45_io_cout)
  );
  FullAdder fa_46 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_46_io_a),
    .io_b(fa_46_io_b),
    .io_cin(fa_46_io_cin),
    .io_sum(fa_46_io_sum),
    .io_cout(fa_46_io_cout)
  );
  FullAdder fa_47 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_47_io_a),
    .io_b(fa_47_io_b),
    .io_cin(fa_47_io_cin),
    .io_sum(fa_47_io_sum),
    .io_cout(fa_47_io_cout)
  );
  FullAdder fa_48 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_48_io_a),
    .io_b(fa_48_io_b),
    .io_cin(fa_48_io_cin),
    .io_sum(fa_48_io_sum),
    .io_cout(fa_48_io_cout)
  );
  FullAdder fa_49 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_49_io_a),
    .io_b(fa_49_io_b),
    .io_cin(fa_49_io_cin),
    .io_sum(fa_49_io_sum),
    .io_cout(fa_49_io_cout)
  );
  FullAdder fa_50 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_50_io_a),
    .io_b(fa_50_io_b),
    .io_cin(fa_50_io_cin),
    .io_sum(fa_50_io_sum),
    .io_cout(fa_50_io_cout)
  );
  FullAdder fa_51 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_51_io_a),
    .io_b(fa_51_io_b),
    .io_cin(fa_51_io_cin),
    .io_sum(fa_51_io_sum),
    .io_cout(fa_51_io_cout)
  );
  FullAdder fa_52 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_52_io_a),
    .io_b(fa_52_io_b),
    .io_cin(fa_52_io_cin),
    .io_sum(fa_52_io_sum),
    .io_cout(fa_52_io_cout)
  );
  FullAdder fa_53 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_53_io_a),
    .io_b(fa_53_io_b),
    .io_cin(fa_53_io_cin),
    .io_sum(fa_53_io_sum),
    .io_cout(fa_53_io_cout)
  );
  FullAdder fa_54 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_54_io_a),
    .io_b(fa_54_io_b),
    .io_cin(fa_54_io_cin),
    .io_sum(fa_54_io_sum),
    .io_cout(fa_54_io_cout)
  );
  FullAdder fa_55 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_55_io_a),
    .io_b(fa_55_io_b),
    .io_cin(fa_55_io_cin),
    .io_sum(fa_55_io_sum),
    .io_cout(fa_55_io_cout)
  );
  FullAdder fa_56 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_56_io_a),
    .io_b(fa_56_io_b),
    .io_cin(fa_56_io_cin),
    .io_sum(fa_56_io_sum),
    .io_cout(fa_56_io_cout)
  );
  FullAdder fa_57 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_57_io_a),
    .io_b(fa_57_io_b),
    .io_cin(fa_57_io_cin),
    .io_sum(fa_57_io_sum),
    .io_cout(fa_57_io_cout)
  );
  FullAdder fa_58 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_58_io_a),
    .io_b(fa_58_io_b),
    .io_cin(fa_58_io_cin),
    .io_sum(fa_58_io_sum),
    .io_cout(fa_58_io_cout)
  );
  FullAdder fa_59 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_59_io_a),
    .io_b(fa_59_io_b),
    .io_cin(fa_59_io_cin),
    .io_sum(fa_59_io_sum),
    .io_cout(fa_59_io_cout)
  );
  FullAdder fa_60 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_60_io_a),
    .io_b(fa_60_io_b),
    .io_cin(fa_60_io_cin),
    .io_sum(fa_60_io_sum),
    .io_cout(fa_60_io_cout)
  );
  FullAdder fa_61 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_61_io_a),
    .io_b(fa_61_io_b),
    .io_cin(fa_61_io_cin),
    .io_sum(fa_61_io_sum),
    .io_cout(fa_61_io_cout)
  );
  FullAdder fa_62 ( // @[src/main/scala/dadda_tree_mult.scala 49:20]
    .io_a(fa_62_io_a),
    .io_b(fa_62_io_b),
    .io_cin(fa_62_io_cin),
    .io_sum(fa_62_io_sum),
    .io_cout(fa_62_io_cout)
  );
  assign io_sum = {io_sum_hi,io_sum_lo}; // @[src/main/scala/dadda_tree_mult.scala 59:21]
  assign io_cout = fa_62_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_io_a = io_a[0]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_io_b = io_b[0]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_io_cin = 1'h0; // @[src/main/scala/dadda_tree_mult.scala 41:21 42:14]
  assign fa_1_io_a = io_a[1]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_1_io_b = io_b[1]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_1_io_cin = fa_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_2_io_a = io_a[2]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_2_io_b = io_b[2]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_2_io_cin = fa_1_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_3_io_a = io_a[3]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_3_io_b = io_b[3]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_3_io_cin = fa_2_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_4_io_a = io_a[4]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_4_io_b = io_b[4]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_4_io_cin = fa_3_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_5_io_a = io_a[5]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_5_io_b = io_b[5]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_5_io_cin = fa_4_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_6_io_a = io_a[6]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_6_io_b = io_b[6]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_6_io_cin = fa_5_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_7_io_a = io_a[7]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_7_io_b = io_b[7]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_7_io_cin = fa_6_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_8_io_a = io_a[8]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_8_io_b = io_b[8]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_8_io_cin = fa_7_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_9_io_a = io_a[9]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_9_io_b = io_b[9]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_9_io_cin = fa_8_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_10_io_a = io_a[10]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_10_io_b = io_b[10]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_10_io_cin = fa_9_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_11_io_a = io_a[11]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_11_io_b = io_b[11]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_11_io_cin = fa_10_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_12_io_a = io_a[12]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_12_io_b = io_b[12]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_12_io_cin = fa_11_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_13_io_a = io_a[13]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_13_io_b = io_b[13]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_13_io_cin = fa_12_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_14_io_a = io_a[14]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_14_io_b = io_b[14]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_14_io_cin = fa_13_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_15_io_a = io_a[15]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_15_io_b = io_b[15]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_15_io_cin = fa_14_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_16_io_a = io_a[16]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_16_io_b = io_b[16]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_16_io_cin = fa_15_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_17_io_a = io_a[17]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_17_io_b = io_b[17]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_17_io_cin = fa_16_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_18_io_a = io_a[18]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_18_io_b = io_b[18]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_18_io_cin = fa_17_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_19_io_a = io_a[19]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_19_io_b = io_b[19]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_19_io_cin = fa_18_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_20_io_a = io_a[20]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_20_io_b = io_b[20]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_20_io_cin = fa_19_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_21_io_a = io_a[21]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_21_io_b = io_b[21]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_21_io_cin = fa_20_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_22_io_a = io_a[22]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_22_io_b = io_b[22]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_22_io_cin = fa_21_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_23_io_a = io_a[23]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_23_io_b = io_b[23]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_23_io_cin = fa_22_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_24_io_a = io_a[24]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_24_io_b = io_b[24]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_24_io_cin = fa_23_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_25_io_a = io_a[25]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_25_io_b = io_b[25]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_25_io_cin = fa_24_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_26_io_a = io_a[26]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_26_io_b = io_b[26]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_26_io_cin = fa_25_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_27_io_a = io_a[27]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_27_io_b = io_b[27]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_27_io_cin = fa_26_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_28_io_a = io_a[28]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_28_io_b = io_b[28]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_28_io_cin = fa_27_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_29_io_a = io_a[29]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_29_io_b = io_b[29]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_29_io_cin = fa_28_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_30_io_a = io_a[30]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_30_io_b = io_b[30]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_30_io_cin = fa_29_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_31_io_a = io_a[31]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_31_io_b = io_b[31]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_31_io_cin = fa_30_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_32_io_a = io_a[32]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_32_io_b = io_b[32]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_32_io_cin = fa_31_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_33_io_a = io_a[33]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_33_io_b = io_b[33]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_33_io_cin = fa_32_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_34_io_a = io_a[34]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_34_io_b = io_b[34]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_34_io_cin = fa_33_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_35_io_a = io_a[35]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_35_io_b = io_b[35]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_35_io_cin = fa_34_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_36_io_a = io_a[36]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_36_io_b = io_b[36]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_36_io_cin = fa_35_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_37_io_a = io_a[37]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_37_io_b = io_b[37]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_37_io_cin = fa_36_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_38_io_a = io_a[38]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_38_io_b = io_b[38]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_38_io_cin = fa_37_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_39_io_a = io_a[39]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_39_io_b = io_b[39]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_39_io_cin = fa_38_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_40_io_a = io_a[40]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_40_io_b = io_b[40]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_40_io_cin = fa_39_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_41_io_a = io_a[41]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_41_io_b = io_b[41]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_41_io_cin = fa_40_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_42_io_a = io_a[42]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_42_io_b = io_b[42]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_42_io_cin = fa_41_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_43_io_a = io_a[43]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_43_io_b = io_b[43]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_43_io_cin = fa_42_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_44_io_a = io_a[44]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_44_io_b = io_b[44]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_44_io_cin = fa_43_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_45_io_a = io_a[45]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_45_io_b = io_b[45]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_45_io_cin = fa_44_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_46_io_a = io_a[46]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_46_io_b = io_b[46]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_46_io_cin = fa_45_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_47_io_a = io_a[47]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_47_io_b = io_b[47]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_47_io_cin = fa_46_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_48_io_a = io_a[48]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_48_io_b = io_b[48]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_48_io_cin = fa_47_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_49_io_a = io_a[49]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_49_io_b = io_b[49]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_49_io_cin = fa_48_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_50_io_a = io_a[50]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_50_io_b = io_b[50]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_50_io_cin = fa_49_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_51_io_a = io_a[51]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_51_io_b = io_b[51]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_51_io_cin = fa_50_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_52_io_a = io_a[52]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_52_io_b = io_b[52]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_52_io_cin = fa_51_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_53_io_a = io_a[53]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_53_io_b = io_b[53]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_53_io_cin = fa_52_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_54_io_a = io_a[54]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_54_io_b = io_b[54]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_54_io_cin = fa_53_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_55_io_a = io_a[55]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_55_io_b = io_b[55]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_55_io_cin = fa_54_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_56_io_a = io_a[56]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_56_io_b = io_b[56]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_56_io_cin = fa_55_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_57_io_a = io_a[57]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_57_io_b = io_b[57]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_57_io_cin = fa_56_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_58_io_a = io_a[58]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_58_io_b = io_b[58]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_58_io_cin = fa_57_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_59_io_a = io_a[59]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_59_io_b = io_b[59]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_59_io_cin = fa_58_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_60_io_a = io_a[60]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_60_io_b = io_b[60]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_60_io_cin = fa_59_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_61_io_a = io_a[61]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_61_io_b = io_b[61]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_61_io_cin = fa_60_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
  assign fa_62_io_a = io_a[62]; // @[src/main/scala/dadda_tree_mult.scala 50:20]
  assign fa_62_io_b = io_b[62]; // @[src/main/scala/dadda_tree_mult.scala 51:20]
  assign fa_62_io_cin = fa_61_io_cout; // @[src/main/scala/dadda_tree_mult.scala 41:21 55:20]
endmodule
module DaddaTreeMultiplier(
  input         clock,
  input         reset,
  input  [31:0] io_a, // @[src/main/scala/dadda_tree_mult.scala 64:15]
  input  [31:0] io_b, // @[src/main/scala/dadda_tree_mult.scala 64:15]
  output [63:0] io_product // @[src/main/scala/dadda_tree_mult.scala 64:15]
);
  wire [62:0] io_product_rca_io_a; // @[src/main/scala/dadda_tree_mult.scala 163:21]
  wire [62:0] io_product_rca_io_b; // @[src/main/scala/dadda_tree_mult.scala 163:21]
  wire [62:0] io_product_rca_io_sum; // @[src/main/scala/dadda_tree_mult.scala 163:21]
  wire  io_product_rca_io_cout; // @[src/main/scala/dadda_tree_mult.scala 163:21]
  wire  partials_x_bool_0 = io_a[0]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_1 = io_a[1]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_2 = io_a[2]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_3 = io_a[3]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_4 = io_a[4]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_5 = io_a[5]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_6 = io_a[6]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_7 = io_a[7]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_8 = io_a[8]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_9 = io_a[9]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_10 = io_a[10]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_11 = io_a[11]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_12 = io_a[12]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_13 = io_a[13]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_14 = io_a[14]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_15 = io_a[15]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_16 = io_a[16]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_17 = io_a[17]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_18 = io_a[18]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_19 = io_a[19]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_20 = io_a[20]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_21 = io_a[21]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_22 = io_a[22]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_23 = io_a[23]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_24 = io_a[24]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_25 = io_a[25]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_26 = io_a[26]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_27 = io_a[27]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_28 = io_a[28]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_29 = io_a[29]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_30 = io_a[30]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_x_bool_31 = io_a[31]; // @[src/main/scala/dadda_tree_mult.scala 93:20]
  wire  partials_y_bool_31 = io_b[0]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_30 = io_b[1]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_29 = io_b[2]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_28 = io_b[3]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_27 = io_b[4]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_26 = io_b[5]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_25 = io_b[6]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_24 = io_b[7]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_23 = io_b[8]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_22 = io_b[9]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_21 = io_b[10]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_20 = io_b[11]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_19 = io_b[12]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_18 = io_b[13]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_17 = io_b[14]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_16 = io_b[15]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_15 = io_b[16]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_14 = io_b[17]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_13 = io_b[18]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_12 = io_b[19]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_11 = io_b[20]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_10 = io_b[21]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_9 = io_b[22]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_8 = io_b[23]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_7 = io_b[24]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_6 = io_b[25]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_5 = io_b[26]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_4 = io_b[27]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_3 = io_b[28]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_2 = io_b[29]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_1 = io_b[30]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_y_bool_0 = io_b[31]; // @[src/main/scala/dadda_tree_mult.scala 94:20]
  wire  partials_62_0 = partials_x_bool_31 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_61_0 = partials_x_bool_30 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_61_1 = partials_x_bool_31 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_60_0 = partials_x_bool_29 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_60_1 = partials_x_bool_30 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_60_2 = partials_x_bool_31 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_59_0 = partials_x_bool_28 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_59_1 = partials_x_bool_29 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_59_2 = partials_x_bool_30 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_59_3 = partials_x_bool_31 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_58_0 = partials_x_bool_27 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_58_1 = partials_x_bool_28 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_58_2 = partials_x_bool_29 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_58_3 = partials_x_bool_30 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_58_4 = partials_x_bool_31 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_57_0 = partials_x_bool_26 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_57_1 = partials_x_bool_27 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_57_2 = partials_x_bool_28 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_57_3 = partials_x_bool_29 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_57_4 = partials_x_bool_30 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_57_5 = partials_x_bool_31 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_56_0 = partials_x_bool_25 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_56_1 = partials_x_bool_26 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_56_2 = partials_x_bool_27 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_56_3 = partials_x_bool_28 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_56_4 = partials_x_bool_29 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_56_5 = partials_x_bool_30 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_56_6 = partials_x_bool_31 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_55_0 = partials_x_bool_24 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_55_1 = partials_x_bool_25 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_55_2 = partials_x_bool_26 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_55_3 = partials_x_bool_27 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_55_4 = partials_x_bool_28 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_55_5 = partials_x_bool_29 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_55_6 = partials_x_bool_30 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_55_7 = partials_x_bool_31 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_54_0 = partials_x_bool_23 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_54_1 = partials_x_bool_24 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_54_2 = partials_x_bool_25 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_54_3 = partials_x_bool_26 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_54_4 = partials_x_bool_27 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_54_5 = partials_x_bool_28 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_54_6 = partials_x_bool_29 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_54_7 = partials_x_bool_30 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_54_8 = partials_x_bool_31 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_0 = partials_x_bool_22 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_1 = partials_x_bool_23 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_2 = partials_x_bool_24 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_3 = partials_x_bool_25 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_4 = partials_x_bool_26 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_5 = partials_x_bool_27 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_6 = partials_x_bool_28 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_7 = partials_x_bool_29 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_8 = partials_x_bool_30 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_53_9 = partials_x_bool_31 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_0 = partials_x_bool_21 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_1 = partials_x_bool_22 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_2 = partials_x_bool_23 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_3 = partials_x_bool_24 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_4 = partials_x_bool_25 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_5 = partials_x_bool_26 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_6 = partials_x_bool_27 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_7 = partials_x_bool_28 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_8 = partials_x_bool_29 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_9 = partials_x_bool_30 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_52_10 = partials_x_bool_31 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_0 = partials_x_bool_20 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_1 = partials_x_bool_21 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_2 = partials_x_bool_22 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_3 = partials_x_bool_23 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_4 = partials_x_bool_24 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_5 = partials_x_bool_25 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_6 = partials_x_bool_26 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_7 = partials_x_bool_27 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_8 = partials_x_bool_28 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_9 = partials_x_bool_29 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_10 = partials_x_bool_30 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_51_11 = partials_x_bool_31 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_0 = partials_x_bool_19 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_1 = partials_x_bool_20 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_2 = partials_x_bool_21 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_3 = partials_x_bool_22 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_4 = partials_x_bool_23 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_5 = partials_x_bool_24 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_6 = partials_x_bool_25 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_7 = partials_x_bool_26 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_8 = partials_x_bool_27 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_9 = partials_x_bool_28 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_10 = partials_x_bool_29 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_11 = partials_x_bool_30 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_50_12 = partials_x_bool_31 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_0 = partials_x_bool_18 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_1 = partials_x_bool_19 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_2 = partials_x_bool_20 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_3 = partials_x_bool_21 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_4 = partials_x_bool_22 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_5 = partials_x_bool_23 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_6 = partials_x_bool_24 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_7 = partials_x_bool_25 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_8 = partials_x_bool_26 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_9 = partials_x_bool_27 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_10 = partials_x_bool_28 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_11 = partials_x_bool_29 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_12 = partials_x_bool_30 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_49_13 = partials_x_bool_31 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_0 = partials_x_bool_17 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_1 = partials_x_bool_18 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_2 = partials_x_bool_19 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_3 = partials_x_bool_20 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_4 = partials_x_bool_21 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_5 = partials_x_bool_22 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_6 = partials_x_bool_23 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_7 = partials_x_bool_24 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_8 = partials_x_bool_25 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_9 = partials_x_bool_26 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_10 = partials_x_bool_27 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_11 = partials_x_bool_28 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_12 = partials_x_bool_29 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_13 = partials_x_bool_30 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_48_14 = partials_x_bool_31 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_0 = partials_x_bool_16 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_1 = partials_x_bool_17 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_2 = partials_x_bool_18 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_3 = partials_x_bool_19 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_4 = partials_x_bool_20 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_5 = partials_x_bool_21 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_6 = partials_x_bool_22 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_7 = partials_x_bool_23 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_8 = partials_x_bool_24 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_9 = partials_x_bool_25 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_10 = partials_x_bool_26 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_11 = partials_x_bool_27 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_12 = partials_x_bool_28 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_13 = partials_x_bool_29 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_14 = partials_x_bool_30 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_47_15 = partials_x_bool_31 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_0 = partials_x_bool_15 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_1 = partials_x_bool_16 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_2 = partials_x_bool_17 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_3 = partials_x_bool_18 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_4 = partials_x_bool_19 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_5 = partials_x_bool_20 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_6 = partials_x_bool_21 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_7 = partials_x_bool_22 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_8 = partials_x_bool_23 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_9 = partials_x_bool_24 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_10 = partials_x_bool_25 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_11 = partials_x_bool_26 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_12 = partials_x_bool_27 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_13 = partials_x_bool_28 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_14 = partials_x_bool_29 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_15 = partials_x_bool_30 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_46_16 = partials_x_bool_31 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_0 = partials_x_bool_14 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_1 = partials_x_bool_15 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_2 = partials_x_bool_16 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_3 = partials_x_bool_17 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_4 = partials_x_bool_18 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_5 = partials_x_bool_19 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_6 = partials_x_bool_20 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_7 = partials_x_bool_21 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_8 = partials_x_bool_22 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_9 = partials_x_bool_23 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_10 = partials_x_bool_24 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_11 = partials_x_bool_25 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_12 = partials_x_bool_26 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_13 = partials_x_bool_27 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_14 = partials_x_bool_28 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_15 = partials_x_bool_29 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_16 = partials_x_bool_30 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_45_17 = partials_x_bool_31 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_0 = partials_x_bool_13 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_1 = partials_x_bool_14 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_2 = partials_x_bool_15 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_3 = partials_x_bool_16 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_4 = partials_x_bool_17 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_5 = partials_x_bool_18 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_6 = partials_x_bool_19 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_7 = partials_x_bool_20 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_8 = partials_x_bool_21 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_9 = partials_x_bool_22 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_10 = partials_x_bool_23 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_11 = partials_x_bool_24 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_12 = partials_x_bool_25 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_13 = partials_x_bool_26 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_14 = partials_x_bool_27 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_15 = partials_x_bool_28 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_16 = partials_x_bool_29 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_17 = partials_x_bool_30 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_44_18 = partials_x_bool_31 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_0 = partials_x_bool_12 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_1 = partials_x_bool_13 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_2 = partials_x_bool_14 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_3 = partials_x_bool_15 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_4 = partials_x_bool_16 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_5 = partials_x_bool_17 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_6 = partials_x_bool_18 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_7 = partials_x_bool_19 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_8 = partials_x_bool_20 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_9 = partials_x_bool_21 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_10 = partials_x_bool_22 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_11 = partials_x_bool_23 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_12 = partials_x_bool_24 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_13 = partials_x_bool_25 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_14 = partials_x_bool_26 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_15 = partials_x_bool_27 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_16 = partials_x_bool_28 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_17 = partials_x_bool_29 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_18 = partials_x_bool_30 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_43_19 = partials_x_bool_31 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_0 = partials_x_bool_11 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_1 = partials_x_bool_12 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_2 = partials_x_bool_13 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_3 = partials_x_bool_14 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_4 = partials_x_bool_15 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_5 = partials_x_bool_16 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_6 = partials_x_bool_17 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_7 = partials_x_bool_18 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_8 = partials_x_bool_19 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_9 = partials_x_bool_20 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_10 = partials_x_bool_21 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_11 = partials_x_bool_22 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_12 = partials_x_bool_23 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_13 = partials_x_bool_24 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_14 = partials_x_bool_25 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_15 = partials_x_bool_26 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_16 = partials_x_bool_27 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_17 = partials_x_bool_28 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_18 = partials_x_bool_29 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_19 = partials_x_bool_30 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_42_20 = partials_x_bool_31 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_0 = partials_x_bool_10 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_1 = partials_x_bool_11 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_2 = partials_x_bool_12 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_3 = partials_x_bool_13 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_4 = partials_x_bool_14 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_5 = partials_x_bool_15 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_6 = partials_x_bool_16 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_7 = partials_x_bool_17 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_8 = partials_x_bool_18 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_9 = partials_x_bool_19 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_10 = partials_x_bool_20 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_11 = partials_x_bool_21 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_12 = partials_x_bool_22 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_13 = partials_x_bool_23 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_14 = partials_x_bool_24 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_15 = partials_x_bool_25 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_16 = partials_x_bool_26 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_17 = partials_x_bool_27 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_18 = partials_x_bool_28 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_19 = partials_x_bool_29 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_20 = partials_x_bool_30 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_41_21 = partials_x_bool_31 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_0 = partials_x_bool_9 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_1 = partials_x_bool_10 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_2 = partials_x_bool_11 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_3 = partials_x_bool_12 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_4 = partials_x_bool_13 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_5 = partials_x_bool_14 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_6 = partials_x_bool_15 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_7 = partials_x_bool_16 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_8 = partials_x_bool_17 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_9 = partials_x_bool_18 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_10 = partials_x_bool_19 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_11 = partials_x_bool_20 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_12 = partials_x_bool_21 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_13 = partials_x_bool_22 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_14 = partials_x_bool_23 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_15 = partials_x_bool_24 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_16 = partials_x_bool_25 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_17 = partials_x_bool_26 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_18 = partials_x_bool_27 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_19 = partials_x_bool_28 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_20 = partials_x_bool_29 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_21 = partials_x_bool_30 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_40_22 = partials_x_bool_31 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_0 = partials_x_bool_8 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_1 = partials_x_bool_9 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_2 = partials_x_bool_10 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_3 = partials_x_bool_11 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_4 = partials_x_bool_12 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_5 = partials_x_bool_13 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_6 = partials_x_bool_14 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_7 = partials_x_bool_15 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_8 = partials_x_bool_16 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_9 = partials_x_bool_17 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_10 = partials_x_bool_18 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_11 = partials_x_bool_19 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_12 = partials_x_bool_20 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_13 = partials_x_bool_21 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_14 = partials_x_bool_22 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_15 = partials_x_bool_23 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_16 = partials_x_bool_24 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_17 = partials_x_bool_25 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_18 = partials_x_bool_26 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_19 = partials_x_bool_27 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_20 = partials_x_bool_28 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_21 = partials_x_bool_29 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_22 = partials_x_bool_30 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_39_23 = partials_x_bool_31 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_0 = partials_x_bool_7 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_1 = partials_x_bool_8 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_2 = partials_x_bool_9 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_3 = partials_x_bool_10 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_4 = partials_x_bool_11 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_5 = partials_x_bool_12 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_6 = partials_x_bool_13 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_7 = partials_x_bool_14 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_8 = partials_x_bool_15 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_9 = partials_x_bool_16 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_10 = partials_x_bool_17 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_11 = partials_x_bool_18 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_12 = partials_x_bool_19 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_13 = partials_x_bool_20 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_14 = partials_x_bool_21 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_15 = partials_x_bool_22 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_16 = partials_x_bool_23 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_17 = partials_x_bool_24 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_18 = partials_x_bool_25 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_19 = partials_x_bool_26 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_20 = partials_x_bool_27 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_21 = partials_x_bool_28 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_22 = partials_x_bool_29 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_23 = partials_x_bool_30 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_38_24 = partials_x_bool_31 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_0 = partials_x_bool_6 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_1 = partials_x_bool_7 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_2 = partials_x_bool_8 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_3 = partials_x_bool_9 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_4 = partials_x_bool_10 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_5 = partials_x_bool_11 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_6 = partials_x_bool_12 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_7 = partials_x_bool_13 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_8 = partials_x_bool_14 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_9 = partials_x_bool_15 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_10 = partials_x_bool_16 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_11 = partials_x_bool_17 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_12 = partials_x_bool_18 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_13 = partials_x_bool_19 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_14 = partials_x_bool_20 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_15 = partials_x_bool_21 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_16 = partials_x_bool_22 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_17 = partials_x_bool_23 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_18 = partials_x_bool_24 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_19 = partials_x_bool_25 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_20 = partials_x_bool_26 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_21 = partials_x_bool_27 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_22 = partials_x_bool_28 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_23 = partials_x_bool_29 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_24 = partials_x_bool_30 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_37_25 = partials_x_bool_31 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_0 = partials_x_bool_5 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_1 = partials_x_bool_6 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_2 = partials_x_bool_7 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_3 = partials_x_bool_8 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_4 = partials_x_bool_9 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_5 = partials_x_bool_10 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_6 = partials_x_bool_11 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_7 = partials_x_bool_12 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_8 = partials_x_bool_13 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_9 = partials_x_bool_14 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_10 = partials_x_bool_15 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_11 = partials_x_bool_16 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_12 = partials_x_bool_17 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_13 = partials_x_bool_18 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_14 = partials_x_bool_19 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_15 = partials_x_bool_20 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_16 = partials_x_bool_21 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_17 = partials_x_bool_22 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_18 = partials_x_bool_23 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_19 = partials_x_bool_24 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_20 = partials_x_bool_25 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_21 = partials_x_bool_26 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_22 = partials_x_bool_27 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_23 = partials_x_bool_28 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_24 = partials_x_bool_29 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_25 = partials_x_bool_30 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_36_26 = partials_x_bool_31 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_0 = partials_x_bool_4 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_1 = partials_x_bool_5 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_2 = partials_x_bool_6 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_3 = partials_x_bool_7 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_4 = partials_x_bool_8 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_5 = partials_x_bool_9 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_6 = partials_x_bool_10 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_7 = partials_x_bool_11 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_8 = partials_x_bool_12 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_9 = partials_x_bool_13 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_10 = partials_x_bool_14 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_11 = partials_x_bool_15 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_12 = partials_x_bool_16 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_13 = partials_x_bool_17 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_14 = partials_x_bool_18 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_15 = partials_x_bool_19 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_16 = partials_x_bool_20 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_17 = partials_x_bool_21 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_18 = partials_x_bool_22 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_19 = partials_x_bool_23 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_20 = partials_x_bool_24 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_21 = partials_x_bool_25 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_22 = partials_x_bool_26 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_23 = partials_x_bool_27 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_24 = partials_x_bool_28 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_25 = partials_x_bool_29 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_26 = partials_x_bool_30 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_35_27 = partials_x_bool_31 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_0 = partials_x_bool_3 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_1 = partials_x_bool_4 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_2 = partials_x_bool_5 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_3 = partials_x_bool_6 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_4 = partials_x_bool_7 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_5 = partials_x_bool_8 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_6 = partials_x_bool_9 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_7 = partials_x_bool_10 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_8 = partials_x_bool_11 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_9 = partials_x_bool_12 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_10 = partials_x_bool_13 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_11 = partials_x_bool_14 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_12 = partials_x_bool_15 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_13 = partials_x_bool_16 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_14 = partials_x_bool_17 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_15 = partials_x_bool_18 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_16 = partials_x_bool_19 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_17 = partials_x_bool_20 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_18 = partials_x_bool_21 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_19 = partials_x_bool_22 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_20 = partials_x_bool_23 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_21 = partials_x_bool_24 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_22 = partials_x_bool_25 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_23 = partials_x_bool_26 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_24 = partials_x_bool_27 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_25 = partials_x_bool_28 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_26 = partials_x_bool_29 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_27 = partials_x_bool_30 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_34_28 = partials_x_bool_31 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_0 = partials_x_bool_2 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_1 = partials_x_bool_3 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_2 = partials_x_bool_4 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_3 = partials_x_bool_5 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_4 = partials_x_bool_6 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_5 = partials_x_bool_7 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_6 = partials_x_bool_8 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_7 = partials_x_bool_9 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_8 = partials_x_bool_10 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_9 = partials_x_bool_11 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_10 = partials_x_bool_12 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_11 = partials_x_bool_13 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_12 = partials_x_bool_14 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_13 = partials_x_bool_15 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_14 = partials_x_bool_16 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_15 = partials_x_bool_17 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_16 = partials_x_bool_18 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_17 = partials_x_bool_19 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_18 = partials_x_bool_20 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_19 = partials_x_bool_21 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_20 = partials_x_bool_22 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_21 = partials_x_bool_23 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_22 = partials_x_bool_24 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_23 = partials_x_bool_25 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_24 = partials_x_bool_26 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_25 = partials_x_bool_27 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_26 = partials_x_bool_28 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_27 = partials_x_bool_29 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_28 = partials_x_bool_30 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_33_29 = partials_x_bool_31 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_0 = partials_x_bool_1 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_1 = partials_x_bool_2 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_2 = partials_x_bool_3 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_3 = partials_x_bool_4 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_4 = partials_x_bool_5 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_5 = partials_x_bool_6 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_6 = partials_x_bool_7 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_7 = partials_x_bool_8 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_8 = partials_x_bool_9 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_9 = partials_x_bool_10 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_10 = partials_x_bool_11 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_11 = partials_x_bool_12 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_12 = partials_x_bool_13 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_13 = partials_x_bool_14 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_14 = partials_x_bool_15 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_15 = partials_x_bool_16 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_16 = partials_x_bool_17 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_17 = partials_x_bool_18 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_18 = partials_x_bool_19 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_19 = partials_x_bool_20 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_20 = partials_x_bool_21 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_21 = partials_x_bool_22 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_22 = partials_x_bool_23 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_23 = partials_x_bool_24 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_24 = partials_x_bool_25 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_25 = partials_x_bool_26 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_26 = partials_x_bool_27 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_27 = partials_x_bool_28 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_28 = partials_x_bool_29 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_29 = partials_x_bool_30 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_32_30 = partials_x_bool_31 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_0 = partials_x_bool_0 & partials_y_bool_0; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_1 = partials_x_bool_1 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_2 = partials_x_bool_2 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_3 = partials_x_bool_3 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_4 = partials_x_bool_4 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_5 = partials_x_bool_5 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_6 = partials_x_bool_6 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_7 = partials_x_bool_7 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_8 = partials_x_bool_8 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_9 = partials_x_bool_9 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_10 = partials_x_bool_10 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_11 = partials_x_bool_11 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_12 = partials_x_bool_12 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_13 = partials_x_bool_13 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_14 = partials_x_bool_14 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_15 = partials_x_bool_15 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_16 = partials_x_bool_16 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_17 = partials_x_bool_17 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_18 = partials_x_bool_18 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_19 = partials_x_bool_19 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_20 = partials_x_bool_20 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_21 = partials_x_bool_21 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_22 = partials_x_bool_22 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_23 = partials_x_bool_23 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_24 = partials_x_bool_24 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_25 = partials_x_bool_25 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_26 = partials_x_bool_26 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_27 = partials_x_bool_27 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_28 = partials_x_bool_28 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_29 = partials_x_bool_29 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_30 = partials_x_bool_30 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_31_31 = partials_x_bool_31 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 96:112]
  wire  partials_30_0 = partials_x_bool_0 & partials_y_bool_1; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_1 = partials_x_bool_1 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_2 = partials_x_bool_2 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_3 = partials_x_bool_3 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_4 = partials_x_bool_4 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_5 = partials_x_bool_5 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_6 = partials_x_bool_6 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_7 = partials_x_bool_7 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_8 = partials_x_bool_8 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_9 = partials_x_bool_9 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_10 = partials_x_bool_10 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_11 = partials_x_bool_11 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_12 = partials_x_bool_12 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_13 = partials_x_bool_13 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_14 = partials_x_bool_14 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_15 = partials_x_bool_15 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_16 = partials_x_bool_16 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_17 = partials_x_bool_17 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_18 = partials_x_bool_18 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_19 = partials_x_bool_19 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_20 = partials_x_bool_20 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_21 = partials_x_bool_21 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_22 = partials_x_bool_22 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_23 = partials_x_bool_23 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_24 = partials_x_bool_24 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_25 = partials_x_bool_25 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_26 = partials_x_bool_26 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_27 = partials_x_bool_27 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_28 = partials_x_bool_28 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_29 = partials_x_bool_29 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_30_30 = partials_x_bool_30 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_0 = partials_x_bool_0 & partials_y_bool_2; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_1 = partials_x_bool_1 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_2 = partials_x_bool_2 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_3 = partials_x_bool_3 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_4 = partials_x_bool_4 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_5 = partials_x_bool_5 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_6 = partials_x_bool_6 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_7 = partials_x_bool_7 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_8 = partials_x_bool_8 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_9 = partials_x_bool_9 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_10 = partials_x_bool_10 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_11 = partials_x_bool_11 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_12 = partials_x_bool_12 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_13 = partials_x_bool_13 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_14 = partials_x_bool_14 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_15 = partials_x_bool_15 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_16 = partials_x_bool_16 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_17 = partials_x_bool_17 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_18 = partials_x_bool_18 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_19 = partials_x_bool_19 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_20 = partials_x_bool_20 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_21 = partials_x_bool_21 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_22 = partials_x_bool_22 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_23 = partials_x_bool_23 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_24 = partials_x_bool_24 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_25 = partials_x_bool_25 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_26 = partials_x_bool_26 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_27 = partials_x_bool_27 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_28 = partials_x_bool_28 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_29_29 = partials_x_bool_29 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_0 = partials_x_bool_0 & partials_y_bool_3; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_1 = partials_x_bool_1 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_2 = partials_x_bool_2 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_3 = partials_x_bool_3 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_4 = partials_x_bool_4 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_5 = partials_x_bool_5 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_6 = partials_x_bool_6 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_7 = partials_x_bool_7 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_8 = partials_x_bool_8 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_9 = partials_x_bool_9 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_10 = partials_x_bool_10 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_11 = partials_x_bool_11 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_12 = partials_x_bool_12 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_13 = partials_x_bool_13 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_14 = partials_x_bool_14 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_15 = partials_x_bool_15 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_16 = partials_x_bool_16 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_17 = partials_x_bool_17 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_18 = partials_x_bool_18 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_19 = partials_x_bool_19 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_20 = partials_x_bool_20 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_21 = partials_x_bool_21 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_22 = partials_x_bool_22 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_23 = partials_x_bool_23 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_24 = partials_x_bool_24 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_25 = partials_x_bool_25 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_26 = partials_x_bool_26 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_27 = partials_x_bool_27 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_28_28 = partials_x_bool_28 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_0 = partials_x_bool_0 & partials_y_bool_4; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_1 = partials_x_bool_1 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_2 = partials_x_bool_2 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_3 = partials_x_bool_3 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_4 = partials_x_bool_4 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_5 = partials_x_bool_5 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_6 = partials_x_bool_6 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_7 = partials_x_bool_7 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_8 = partials_x_bool_8 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_9 = partials_x_bool_9 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_10 = partials_x_bool_10 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_11 = partials_x_bool_11 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_12 = partials_x_bool_12 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_13 = partials_x_bool_13 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_14 = partials_x_bool_14 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_15 = partials_x_bool_15 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_16 = partials_x_bool_16 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_17 = partials_x_bool_17 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_18 = partials_x_bool_18 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_19 = partials_x_bool_19 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_20 = partials_x_bool_20 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_21 = partials_x_bool_21 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_22 = partials_x_bool_22 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_23 = partials_x_bool_23 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_24 = partials_x_bool_24 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_25 = partials_x_bool_25 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_26 = partials_x_bool_26 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_27_27 = partials_x_bool_27 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_0 = partials_x_bool_0 & partials_y_bool_5; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_1 = partials_x_bool_1 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_2 = partials_x_bool_2 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_3 = partials_x_bool_3 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_4 = partials_x_bool_4 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_5 = partials_x_bool_5 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_6 = partials_x_bool_6 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_7 = partials_x_bool_7 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_8 = partials_x_bool_8 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_9 = partials_x_bool_9 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_10 = partials_x_bool_10 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_11 = partials_x_bool_11 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_12 = partials_x_bool_12 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_13 = partials_x_bool_13 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_14 = partials_x_bool_14 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_15 = partials_x_bool_15 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_16 = partials_x_bool_16 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_17 = partials_x_bool_17 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_18 = partials_x_bool_18 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_19 = partials_x_bool_19 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_20 = partials_x_bool_20 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_21 = partials_x_bool_21 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_22 = partials_x_bool_22 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_23 = partials_x_bool_23 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_24 = partials_x_bool_24 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_25 = partials_x_bool_25 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_26_26 = partials_x_bool_26 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_0 = partials_x_bool_0 & partials_y_bool_6; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_1 = partials_x_bool_1 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_2 = partials_x_bool_2 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_3 = partials_x_bool_3 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_4 = partials_x_bool_4 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_5 = partials_x_bool_5 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_6 = partials_x_bool_6 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_7 = partials_x_bool_7 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_8 = partials_x_bool_8 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_9 = partials_x_bool_9 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_10 = partials_x_bool_10 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_11 = partials_x_bool_11 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_12 = partials_x_bool_12 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_13 = partials_x_bool_13 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_14 = partials_x_bool_14 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_15 = partials_x_bool_15 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_16 = partials_x_bool_16 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_17 = partials_x_bool_17 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_18 = partials_x_bool_18 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_19 = partials_x_bool_19 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_20 = partials_x_bool_20 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_21 = partials_x_bool_21 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_22 = partials_x_bool_22 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_23 = partials_x_bool_23 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_24 = partials_x_bool_24 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_25_25 = partials_x_bool_25 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_0 = partials_x_bool_0 & partials_y_bool_7; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_1 = partials_x_bool_1 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_2 = partials_x_bool_2 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_3 = partials_x_bool_3 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_4 = partials_x_bool_4 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_5 = partials_x_bool_5 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_6 = partials_x_bool_6 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_7 = partials_x_bool_7 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_8 = partials_x_bool_8 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_9 = partials_x_bool_9 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_10 = partials_x_bool_10 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_11 = partials_x_bool_11 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_12 = partials_x_bool_12 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_13 = partials_x_bool_13 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_14 = partials_x_bool_14 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_15 = partials_x_bool_15 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_16 = partials_x_bool_16 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_17 = partials_x_bool_17 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_18 = partials_x_bool_18 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_19 = partials_x_bool_19 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_20 = partials_x_bool_20 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_21 = partials_x_bool_21 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_22 = partials_x_bool_22 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_23 = partials_x_bool_23 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_24_24 = partials_x_bool_24 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_0 = partials_x_bool_0 & partials_y_bool_8; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_1 = partials_x_bool_1 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_2 = partials_x_bool_2 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_3 = partials_x_bool_3 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_4 = partials_x_bool_4 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_5 = partials_x_bool_5 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_6 = partials_x_bool_6 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_7 = partials_x_bool_7 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_8 = partials_x_bool_8 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_9 = partials_x_bool_9 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_10 = partials_x_bool_10 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_11 = partials_x_bool_11 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_12 = partials_x_bool_12 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_13 = partials_x_bool_13 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_14 = partials_x_bool_14 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_15 = partials_x_bool_15 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_16 = partials_x_bool_16 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_17 = partials_x_bool_17 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_18 = partials_x_bool_18 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_19 = partials_x_bool_19 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_20 = partials_x_bool_20 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_21 = partials_x_bool_21 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_22 = partials_x_bool_22 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_23_23 = partials_x_bool_23 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_0 = partials_x_bool_0 & partials_y_bool_9; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_1 = partials_x_bool_1 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_2 = partials_x_bool_2 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_3 = partials_x_bool_3 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_4 = partials_x_bool_4 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_5 = partials_x_bool_5 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_6 = partials_x_bool_6 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_7 = partials_x_bool_7 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_8 = partials_x_bool_8 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_9 = partials_x_bool_9 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_10 = partials_x_bool_10 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_11 = partials_x_bool_11 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_12 = partials_x_bool_12 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_13 = partials_x_bool_13 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_14 = partials_x_bool_14 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_15 = partials_x_bool_15 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_16 = partials_x_bool_16 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_17 = partials_x_bool_17 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_18 = partials_x_bool_18 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_19 = partials_x_bool_19 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_20 = partials_x_bool_20 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_21 = partials_x_bool_21 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_22_22 = partials_x_bool_22 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_0 = partials_x_bool_0 & partials_y_bool_10; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_1 = partials_x_bool_1 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_2 = partials_x_bool_2 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_3 = partials_x_bool_3 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_4 = partials_x_bool_4 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_5 = partials_x_bool_5 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_6 = partials_x_bool_6 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_7 = partials_x_bool_7 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_8 = partials_x_bool_8 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_9 = partials_x_bool_9 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_10 = partials_x_bool_10 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_11 = partials_x_bool_11 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_12 = partials_x_bool_12 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_13 = partials_x_bool_13 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_14 = partials_x_bool_14 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_15 = partials_x_bool_15 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_16 = partials_x_bool_16 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_17 = partials_x_bool_17 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_18 = partials_x_bool_18 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_19 = partials_x_bool_19 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_20 = partials_x_bool_20 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_21_21 = partials_x_bool_21 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_0 = partials_x_bool_0 & partials_y_bool_11; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_1 = partials_x_bool_1 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_2 = partials_x_bool_2 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_3 = partials_x_bool_3 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_4 = partials_x_bool_4 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_5 = partials_x_bool_5 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_6 = partials_x_bool_6 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_7 = partials_x_bool_7 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_8 = partials_x_bool_8 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_9 = partials_x_bool_9 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_10 = partials_x_bool_10 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_11 = partials_x_bool_11 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_12 = partials_x_bool_12 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_13 = partials_x_bool_13 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_14 = partials_x_bool_14 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_15 = partials_x_bool_15 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_16 = partials_x_bool_16 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_17 = partials_x_bool_17 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_18 = partials_x_bool_18 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_19 = partials_x_bool_19 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_20_20 = partials_x_bool_20 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_0 = partials_x_bool_0 & partials_y_bool_12; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_1 = partials_x_bool_1 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_2 = partials_x_bool_2 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_3 = partials_x_bool_3 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_4 = partials_x_bool_4 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_5 = partials_x_bool_5 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_6 = partials_x_bool_6 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_7 = partials_x_bool_7 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_8 = partials_x_bool_8 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_9 = partials_x_bool_9 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_10 = partials_x_bool_10 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_11 = partials_x_bool_11 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_12 = partials_x_bool_12 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_13 = partials_x_bool_13 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_14 = partials_x_bool_14 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_15 = partials_x_bool_15 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_16 = partials_x_bool_16 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_17 = partials_x_bool_17 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_18 = partials_x_bool_18 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_19_19 = partials_x_bool_19 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_0 = partials_x_bool_0 & partials_y_bool_13; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_1 = partials_x_bool_1 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_2 = partials_x_bool_2 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_3 = partials_x_bool_3 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_4 = partials_x_bool_4 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_5 = partials_x_bool_5 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_6 = partials_x_bool_6 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_7 = partials_x_bool_7 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_8 = partials_x_bool_8 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_9 = partials_x_bool_9 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_10 = partials_x_bool_10 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_11 = partials_x_bool_11 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_12 = partials_x_bool_12 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_13 = partials_x_bool_13 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_14 = partials_x_bool_14 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_15 = partials_x_bool_15 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_16 = partials_x_bool_16 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_17 = partials_x_bool_17 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_18_18 = partials_x_bool_18 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_0 = partials_x_bool_0 & partials_y_bool_14; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_1 = partials_x_bool_1 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_2 = partials_x_bool_2 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_3 = partials_x_bool_3 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_4 = partials_x_bool_4 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_5 = partials_x_bool_5 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_6 = partials_x_bool_6 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_7 = partials_x_bool_7 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_8 = partials_x_bool_8 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_9 = partials_x_bool_9 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_10 = partials_x_bool_10 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_11 = partials_x_bool_11 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_12 = partials_x_bool_12 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_13 = partials_x_bool_13 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_14 = partials_x_bool_14 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_15 = partials_x_bool_15 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_16 = partials_x_bool_16 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_17_17 = partials_x_bool_17 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_0 = partials_x_bool_0 & partials_y_bool_15; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_1 = partials_x_bool_1 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_2 = partials_x_bool_2 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_3 = partials_x_bool_3 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_4 = partials_x_bool_4 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_5 = partials_x_bool_5 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_6 = partials_x_bool_6 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_7 = partials_x_bool_7 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_8 = partials_x_bool_8 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_9 = partials_x_bool_9 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_10 = partials_x_bool_10 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_11 = partials_x_bool_11 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_12 = partials_x_bool_12 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_13 = partials_x_bool_13 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_14 = partials_x_bool_14 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_15 = partials_x_bool_15 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_16_16 = partials_x_bool_16 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_0 = partials_x_bool_0 & partials_y_bool_16; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_1 = partials_x_bool_1 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_2 = partials_x_bool_2 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_3 = partials_x_bool_3 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_4 = partials_x_bool_4 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_5 = partials_x_bool_5 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_6 = partials_x_bool_6 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_7 = partials_x_bool_7 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_8 = partials_x_bool_8 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_9 = partials_x_bool_9 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_10 = partials_x_bool_10 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_11 = partials_x_bool_11 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_12 = partials_x_bool_12 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_13 = partials_x_bool_13 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_14 = partials_x_bool_14 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_15_15 = partials_x_bool_15 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_0 = partials_x_bool_0 & partials_y_bool_17; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_1 = partials_x_bool_1 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_2 = partials_x_bool_2 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_3 = partials_x_bool_3 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_4 = partials_x_bool_4 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_5 = partials_x_bool_5 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_6 = partials_x_bool_6 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_7 = partials_x_bool_7 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_8 = partials_x_bool_8 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_9 = partials_x_bool_9 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_10 = partials_x_bool_10 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_11 = partials_x_bool_11 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_12 = partials_x_bool_12 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_13 = partials_x_bool_13 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_14_14 = partials_x_bool_14 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_0 = partials_x_bool_0 & partials_y_bool_18; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_1 = partials_x_bool_1 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_2 = partials_x_bool_2 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_3 = partials_x_bool_3 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_4 = partials_x_bool_4 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_5 = partials_x_bool_5 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_6 = partials_x_bool_6 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_7 = partials_x_bool_7 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_8 = partials_x_bool_8 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_9 = partials_x_bool_9 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_10 = partials_x_bool_10 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_11 = partials_x_bool_11 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_12 = partials_x_bool_12 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_13_13 = partials_x_bool_13 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_0 = partials_x_bool_0 & partials_y_bool_19; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_1 = partials_x_bool_1 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_2 = partials_x_bool_2 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_3 = partials_x_bool_3 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_4 = partials_x_bool_4 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_5 = partials_x_bool_5 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_6 = partials_x_bool_6 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_7 = partials_x_bool_7 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_8 = partials_x_bool_8 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_9 = partials_x_bool_9 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_10 = partials_x_bool_10 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_11 = partials_x_bool_11 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_12_12 = partials_x_bool_12 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_0 = partials_x_bool_0 & partials_y_bool_20; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_1 = partials_x_bool_1 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_2 = partials_x_bool_2 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_3 = partials_x_bool_3 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_4 = partials_x_bool_4 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_5 = partials_x_bool_5 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_6 = partials_x_bool_6 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_7 = partials_x_bool_7 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_8 = partials_x_bool_8 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_9 = partials_x_bool_9 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_10 = partials_x_bool_10 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_11_11 = partials_x_bool_11 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_0 = partials_x_bool_0 & partials_y_bool_21; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_1 = partials_x_bool_1 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_2 = partials_x_bool_2 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_3 = partials_x_bool_3 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_4 = partials_x_bool_4 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_5 = partials_x_bool_5 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_6 = partials_x_bool_6 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_7 = partials_x_bool_7 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_8 = partials_x_bool_8 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_9 = partials_x_bool_9 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_10_10 = partials_x_bool_10 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_0 = partials_x_bool_0 & partials_y_bool_22; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_1 = partials_x_bool_1 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_2 = partials_x_bool_2 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_3 = partials_x_bool_3 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_4 = partials_x_bool_4 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_5 = partials_x_bool_5 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_6 = partials_x_bool_6 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_7 = partials_x_bool_7 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_8 = partials_x_bool_8 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_9_9 = partials_x_bool_9 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_8_0 = partials_x_bool_0 & partials_y_bool_23; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_8_1 = partials_x_bool_1 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_8_2 = partials_x_bool_2 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_8_3 = partials_x_bool_3 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_8_4 = partials_x_bool_4 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_8_5 = partials_x_bool_5 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_8_6 = partials_x_bool_6 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_8_7 = partials_x_bool_7 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_8_8 = partials_x_bool_8 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_7_0 = partials_x_bool_0 & partials_y_bool_24; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_7_1 = partials_x_bool_1 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_7_2 = partials_x_bool_2 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_7_3 = partials_x_bool_3 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_7_4 = partials_x_bool_4 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_7_5 = partials_x_bool_5 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_7_6 = partials_x_bool_6 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_7_7 = partials_x_bool_7 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_6_0 = partials_x_bool_0 & partials_y_bool_25; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_6_1 = partials_x_bool_1 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_6_2 = partials_x_bool_2 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_6_3 = partials_x_bool_3 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_6_4 = partials_x_bool_4 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_6_5 = partials_x_bool_5 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_6_6 = partials_x_bool_6 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_5_0 = partials_x_bool_0 & partials_y_bool_26; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_5_1 = partials_x_bool_1 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_5_2 = partials_x_bool_2 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_5_3 = partials_x_bool_3 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_5_4 = partials_x_bool_4 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_5_5 = partials_x_bool_5 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_4_0 = partials_x_bool_0 & partials_y_bool_27; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_4_1 = partials_x_bool_1 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_4_2 = partials_x_bool_2 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_4_3 = partials_x_bool_3 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_4_4 = partials_x_bool_4 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_3_0 = partials_x_bool_0 & partials_y_bool_28; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_3_1 = partials_x_bool_1 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_3_2 = partials_x_bool_2 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_3_3 = partials_x_bool_3 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_2_0 = partials_x_bool_0 & partials_y_bool_29; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_2_1 = partials_x_bool_1 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_2_2 = partials_x_bool_2 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_1_0 = partials_x_bool_0 & partials_y_bool_30; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_1_1 = partials_x_bool_1 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  partials_0_0 = partials_x_bool_0 & partials_y_bool_31; // @[src/main/scala/dadda_tree_mult.scala 97:113]
  wire  reducedPartials_reducedPartials_28_0 = partials_28_0 ^ partials_28_1; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry = partials_28_0 & partials_28_1; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum = reducedPartials_reducedPartials_carry ^ partials_29_0 ^ partials_29_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_1 = reducedPartials_reducedPartials_carry & partials_29_0 | partials_29_0
     & partials_29_1 | reducedPartials_reducedPartials_carry & partials_29_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_29_0 = reducedPartials_reducedPartials_sum ^ partials_29_2; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_2 = reducedPartials_reducedPartials_sum & partials_29_2; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_1 = reducedPartials_reducedPartials_carry_2 ^
    reducedPartials_reducedPartials_carry_1 ^ partials_30_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_3 = reducedPartials_reducedPartials_carry_2 &
    reducedPartials_reducedPartials_carry_1 | reducedPartials_reducedPartials_carry_1 & partials_30_0 |
    reducedPartials_reducedPartials_carry_2 & partials_30_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_2 = reducedPartials_reducedPartials_sum_1 ^ partials_30_1 ^ partials_30_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_4 = reducedPartials_reducedPartials_sum_1 & partials_30_1 | partials_30_1
     & partials_30_2 | reducedPartials_reducedPartials_sum_1 & partials_30_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_30_0 = reducedPartials_reducedPartials_sum_2 ^ partials_30_3; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_5 = reducedPartials_reducedPartials_sum_2 & partials_30_3; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_3 = reducedPartials_reducedPartials_carry_5 ^
    reducedPartials_reducedPartials_carry_4 ^ reducedPartials_reducedPartials_carry_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_6 = reducedPartials_reducedPartials_carry_5 &
    reducedPartials_reducedPartials_carry_4 | reducedPartials_reducedPartials_carry_4 &
    reducedPartials_reducedPartials_carry_3 | reducedPartials_reducedPartials_carry_5 &
    reducedPartials_reducedPartials_carry_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_4 = reducedPartials_reducedPartials_sum_3 ^ partials_31_0 ^ partials_31_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_7 = reducedPartials_reducedPartials_sum_3 & partials_31_0 | partials_31_0
     & partials_31_1 | reducedPartials_reducedPartials_sum_3 & partials_31_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_5 = reducedPartials_reducedPartials_sum_4 ^ partials_31_2 ^ partials_31_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_8 = reducedPartials_reducedPartials_sum_4 & partials_31_2 | partials_31_2
     & partials_31_3 | reducedPartials_reducedPartials_sum_4 & partials_31_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_31_0 = reducedPartials_reducedPartials_sum_5 ^ partials_31_4; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_9 = reducedPartials_reducedPartials_sum_5 & partials_31_4; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_6 = reducedPartials_reducedPartials_carry_9 ^
    reducedPartials_reducedPartials_carry_8 ^ reducedPartials_reducedPartials_carry_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_10 = reducedPartials_reducedPartials_carry_9 &
    reducedPartials_reducedPartials_carry_8 | reducedPartials_reducedPartials_carry_8 &
    reducedPartials_reducedPartials_carry_7 | reducedPartials_reducedPartials_carry_9 &
    reducedPartials_reducedPartials_carry_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_7 = reducedPartials_reducedPartials_sum_6 ^
    reducedPartials_reducedPartials_carry_6 ^ partials_32_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_11 = reducedPartials_reducedPartials_sum_6 &
    reducedPartials_reducedPartials_carry_6 | reducedPartials_reducedPartials_carry_6 & partials_32_0 |
    reducedPartials_reducedPartials_sum_6 & partials_32_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_8 = reducedPartials_reducedPartials_sum_7 ^ partials_32_1 ^ partials_32_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_12 = reducedPartials_reducedPartials_sum_7 & partials_32_1 | partials_32_1
     & partials_32_2 | reducedPartials_reducedPartials_sum_7 & partials_32_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_32_0 = reducedPartials_reducedPartials_sum_8 ^ partials_32_3; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_13 = reducedPartials_reducedPartials_sum_8 & partials_32_3; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_9 = reducedPartials_reducedPartials_carry_13 ^
    reducedPartials_reducedPartials_carry_12 ^ reducedPartials_reducedPartials_carry_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_14 = reducedPartials_reducedPartials_carry_13 &
    reducedPartials_reducedPartials_carry_12 | reducedPartials_reducedPartials_carry_12 &
    reducedPartials_reducedPartials_carry_11 | reducedPartials_reducedPartials_carry_13 &
    reducedPartials_reducedPartials_carry_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_10 = reducedPartials_reducedPartials_sum_9 ^
    reducedPartials_reducedPartials_carry_10 ^ partials_33_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_15 = reducedPartials_reducedPartials_sum_9 &
    reducedPartials_reducedPartials_carry_10 | reducedPartials_reducedPartials_carry_10 & partials_33_0 |
    reducedPartials_reducedPartials_sum_9 & partials_33_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_33_0 = reducedPartials_reducedPartials_sum_10 ^ partials_33_1 ^ partials_33_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_16 = reducedPartials_reducedPartials_sum_10 & partials_33_1 |
    partials_33_1 & partials_33_2 | reducedPartials_reducedPartials_sum_10 & partials_33_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_11 = reducedPartials_reducedPartials_carry_16 ^
    reducedPartials_reducedPartials_carry_15 ^ reducedPartials_reducedPartials_carry_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_17 = reducedPartials_reducedPartials_carry_16 &
    reducedPartials_reducedPartials_carry_15 | reducedPartials_reducedPartials_carry_15 &
    reducedPartials_reducedPartials_carry_14 | reducedPartials_reducedPartials_carry_16 &
    reducedPartials_reducedPartials_carry_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_34_0 = reducedPartials_reducedPartials_sum_11 ^ partials_34_0 ^ partials_34_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_18 = reducedPartials_reducedPartials_sum_11 & partials_34_0 |
    partials_34_0 & partials_34_1 | reducedPartials_reducedPartials_sum_11 & partials_34_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_35_0 = reducedPartials_reducedPartials_carry_18 ^
    reducedPartials_reducedPartials_carry_17 ^ partials_35_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_36_0 = reducedPartials_reducedPartials_carry_18 &
    reducedPartials_reducedPartials_carry_17 | reducedPartials_reducedPartials_carry_17 & partials_35_0 |
    reducedPartials_reducedPartials_carry_18 & partials_35_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_19_0 = partials_19_0 ^ partials_19_1; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_19 = partials_19_0 & partials_19_1; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_12 = reducedPartials_reducedPartials_carry_19 ^ partials_20_0 ^
    partials_20_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_20 = reducedPartials_reducedPartials_carry_19 & partials_20_0 |
    partials_20_0 & partials_20_1 | reducedPartials_reducedPartials_carry_19 & partials_20_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_20_0 = reducedPartials_reducedPartials_sum_12 ^ partials_20_2; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_21 = reducedPartials_reducedPartials_sum_12 & partials_20_2; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_13 = reducedPartials_reducedPartials_carry_21 ^
    reducedPartials_reducedPartials_carry_20 ^ partials_21_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_22 = reducedPartials_reducedPartials_carry_21 &
    reducedPartials_reducedPartials_carry_20 | reducedPartials_reducedPartials_carry_20 & partials_21_0 |
    reducedPartials_reducedPartials_carry_21 & partials_21_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_14 = reducedPartials_reducedPartials_sum_13 ^ partials_21_1 ^ partials_21_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_23 = reducedPartials_reducedPartials_sum_13 & partials_21_1 |
    partials_21_1 & partials_21_2 | reducedPartials_reducedPartials_sum_13 & partials_21_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_21_0 = reducedPartials_reducedPartials_sum_14 ^ partials_21_3; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_24 = reducedPartials_reducedPartials_sum_14 & partials_21_3; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_15 = reducedPartials_reducedPartials_carry_24 ^
    reducedPartials_reducedPartials_carry_23 ^ reducedPartials_reducedPartials_carry_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_25 = reducedPartials_reducedPartials_carry_24 &
    reducedPartials_reducedPartials_carry_23 | reducedPartials_reducedPartials_carry_23 &
    reducedPartials_reducedPartials_carry_22 | reducedPartials_reducedPartials_carry_24 &
    reducedPartials_reducedPartials_carry_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_16 = reducedPartials_reducedPartials_sum_15 ^ partials_22_0 ^ partials_22_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_26 = reducedPartials_reducedPartials_sum_15 & partials_22_0 |
    partials_22_0 & partials_22_1 | reducedPartials_reducedPartials_sum_15 & partials_22_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_17 = reducedPartials_reducedPartials_sum_16 ^ partials_22_2 ^ partials_22_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_27 = reducedPartials_reducedPartials_sum_16 & partials_22_2 |
    partials_22_2 & partials_22_3 | reducedPartials_reducedPartials_sum_16 & partials_22_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_22_0 = reducedPartials_reducedPartials_sum_17 ^ partials_22_4; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_28 = reducedPartials_reducedPartials_sum_17 & partials_22_4; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_18 = reducedPartials_reducedPartials_carry_28 ^
    reducedPartials_reducedPartials_carry_27 ^ reducedPartials_reducedPartials_carry_26; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_29 = reducedPartials_reducedPartials_carry_28 &
    reducedPartials_reducedPartials_carry_27 | reducedPartials_reducedPartials_carry_27 &
    reducedPartials_reducedPartials_carry_26 | reducedPartials_reducedPartials_carry_28 &
    reducedPartials_reducedPartials_carry_26; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_19 = reducedPartials_reducedPartials_sum_18 ^
    reducedPartials_reducedPartials_carry_25 ^ partials_23_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_30 = reducedPartials_reducedPartials_sum_18 &
    reducedPartials_reducedPartials_carry_25 | reducedPartials_reducedPartials_carry_25 & partials_23_0 |
    reducedPartials_reducedPartials_sum_18 & partials_23_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_20 = reducedPartials_reducedPartials_sum_19 ^ partials_23_1 ^ partials_23_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_31 = reducedPartials_reducedPartials_sum_19 & partials_23_1 |
    partials_23_1 & partials_23_2 | reducedPartials_reducedPartials_sum_19 & partials_23_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_21 = reducedPartials_reducedPartials_sum_20 ^ partials_23_3 ^ partials_23_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_32 = reducedPartials_reducedPartials_sum_20 & partials_23_3 |
    partials_23_3 & partials_23_4 | reducedPartials_reducedPartials_sum_20 & partials_23_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_23_0 = reducedPartials_reducedPartials_sum_21 ^ partials_23_5; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_33 = reducedPartials_reducedPartials_sum_21 & partials_23_5; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_22 = reducedPartials_reducedPartials_carry_33 ^
    reducedPartials_reducedPartials_carry_32 ^ reducedPartials_reducedPartials_carry_31; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_34 = reducedPartials_reducedPartials_carry_33 &
    reducedPartials_reducedPartials_carry_32 | reducedPartials_reducedPartials_carry_32 &
    reducedPartials_reducedPartials_carry_31 | reducedPartials_reducedPartials_carry_33 &
    reducedPartials_reducedPartials_carry_31; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_23 = reducedPartials_reducedPartials_sum_22 ^
    reducedPartials_reducedPartials_carry_30 ^ reducedPartials_reducedPartials_carry_29; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_35 = reducedPartials_reducedPartials_sum_22 &
    reducedPartials_reducedPartials_carry_30 | reducedPartials_reducedPartials_carry_30 &
    reducedPartials_reducedPartials_carry_29 | reducedPartials_reducedPartials_sum_22 &
    reducedPartials_reducedPartials_carry_29; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_24 = reducedPartials_reducedPartials_sum_23 ^ partials_24_0 ^ partials_24_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_36 = reducedPartials_reducedPartials_sum_23 & partials_24_0 |
    partials_24_0 & partials_24_1 | reducedPartials_reducedPartials_sum_23 & partials_24_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_25 = reducedPartials_reducedPartials_sum_24 ^ partials_24_2 ^ partials_24_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_37 = reducedPartials_reducedPartials_sum_24 & partials_24_2 |
    partials_24_2 & partials_24_3 | reducedPartials_reducedPartials_sum_24 & partials_24_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_26 = reducedPartials_reducedPartials_sum_25 ^ partials_24_4 ^ partials_24_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_38 = reducedPartials_reducedPartials_sum_25 & partials_24_4 |
    partials_24_4 & partials_24_5 | reducedPartials_reducedPartials_sum_25 & partials_24_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_24_0 = reducedPartials_reducedPartials_sum_26 ^ partials_24_6; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_39 = reducedPartials_reducedPartials_sum_26 & partials_24_6; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_27 = reducedPartials_reducedPartials_carry_39 ^
    reducedPartials_reducedPartials_carry_38 ^ reducedPartials_reducedPartials_carry_37; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_40 = reducedPartials_reducedPartials_carry_39 &
    reducedPartials_reducedPartials_carry_38 | reducedPartials_reducedPartials_carry_38 &
    reducedPartials_reducedPartials_carry_37 | reducedPartials_reducedPartials_carry_39 &
    reducedPartials_reducedPartials_carry_37; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_28 = reducedPartials_reducedPartials_sum_27 ^
    reducedPartials_reducedPartials_carry_36 ^ reducedPartials_reducedPartials_carry_35; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_41 = reducedPartials_reducedPartials_sum_27 &
    reducedPartials_reducedPartials_carry_36 | reducedPartials_reducedPartials_carry_36 &
    reducedPartials_reducedPartials_carry_35 | reducedPartials_reducedPartials_sum_27 &
    reducedPartials_reducedPartials_carry_35; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_29 = reducedPartials_reducedPartials_sum_28 ^
    reducedPartials_reducedPartials_carry_34 ^ partials_25_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_42 = reducedPartials_reducedPartials_sum_28 &
    reducedPartials_reducedPartials_carry_34 | reducedPartials_reducedPartials_carry_34 & partials_25_0 |
    reducedPartials_reducedPartials_sum_28 & partials_25_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_30 = reducedPartials_reducedPartials_sum_29 ^ partials_25_1 ^ partials_25_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_43 = reducedPartials_reducedPartials_sum_29 & partials_25_1 |
    partials_25_1 & partials_25_2 | reducedPartials_reducedPartials_sum_29 & partials_25_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_31 = reducedPartials_reducedPartials_sum_30 ^ partials_25_3 ^ partials_25_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_44 = reducedPartials_reducedPartials_sum_30 & partials_25_3 |
    partials_25_3 & partials_25_4 | reducedPartials_reducedPartials_sum_30 & partials_25_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_32 = reducedPartials_reducedPartials_sum_31 ^ partials_25_5 ^ partials_25_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_45 = reducedPartials_reducedPartials_sum_31 & partials_25_5 |
    partials_25_5 & partials_25_6 | reducedPartials_reducedPartials_sum_31 & partials_25_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_25_0 = reducedPartials_reducedPartials_sum_32 ^ partials_25_7; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_46 = reducedPartials_reducedPartials_sum_32 & partials_25_7; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_33 = reducedPartials_reducedPartials_carry_46 ^
    reducedPartials_reducedPartials_carry_45 ^ reducedPartials_reducedPartials_carry_44; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_47 = reducedPartials_reducedPartials_carry_46 &
    reducedPartials_reducedPartials_carry_45 | reducedPartials_reducedPartials_carry_45 &
    reducedPartials_reducedPartials_carry_44 | reducedPartials_reducedPartials_carry_46 &
    reducedPartials_reducedPartials_carry_44; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_34 = reducedPartials_reducedPartials_sum_33 ^
    reducedPartials_reducedPartials_carry_43 ^ reducedPartials_reducedPartials_carry_42; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_48 = reducedPartials_reducedPartials_sum_33 &
    reducedPartials_reducedPartials_carry_43 | reducedPartials_reducedPartials_carry_43 &
    reducedPartials_reducedPartials_carry_42 | reducedPartials_reducedPartials_sum_33 &
    reducedPartials_reducedPartials_carry_42; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_35 = reducedPartials_reducedPartials_sum_34 ^
    reducedPartials_reducedPartials_carry_41 ^ reducedPartials_reducedPartials_carry_40; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_49 = reducedPartials_reducedPartials_sum_34 &
    reducedPartials_reducedPartials_carry_41 | reducedPartials_reducedPartials_carry_41 &
    reducedPartials_reducedPartials_carry_40 | reducedPartials_reducedPartials_sum_34 &
    reducedPartials_reducedPartials_carry_40; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_36 = reducedPartials_reducedPartials_sum_35 ^ partials_26_0 ^ partials_26_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_50 = reducedPartials_reducedPartials_sum_35 & partials_26_0 |
    partials_26_0 & partials_26_1 | reducedPartials_reducedPartials_sum_35 & partials_26_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_37 = reducedPartials_reducedPartials_sum_36 ^ partials_26_2 ^ partials_26_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_51 = reducedPartials_reducedPartials_sum_36 & partials_26_2 |
    partials_26_2 & partials_26_3 | reducedPartials_reducedPartials_sum_36 & partials_26_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_38 = reducedPartials_reducedPartials_sum_37 ^ partials_26_4 ^ partials_26_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_52 = reducedPartials_reducedPartials_sum_37 & partials_26_4 |
    partials_26_4 & partials_26_5 | reducedPartials_reducedPartials_sum_37 & partials_26_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_39 = reducedPartials_reducedPartials_sum_38 ^ partials_26_6 ^ partials_26_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_53 = reducedPartials_reducedPartials_sum_38 & partials_26_6 |
    partials_26_6 & partials_26_7 | reducedPartials_reducedPartials_sum_38 & partials_26_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_26_0 = reducedPartials_reducedPartials_sum_39 ^ partials_26_8; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_54 = reducedPartials_reducedPartials_sum_39 & partials_26_8; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_40 = reducedPartials_reducedPartials_carry_54 ^
    reducedPartials_reducedPartials_carry_53 ^ reducedPartials_reducedPartials_carry_52; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_55 = reducedPartials_reducedPartials_carry_54 &
    reducedPartials_reducedPartials_carry_53 | reducedPartials_reducedPartials_carry_53 &
    reducedPartials_reducedPartials_carry_52 | reducedPartials_reducedPartials_carry_54 &
    reducedPartials_reducedPartials_carry_52; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_41 = reducedPartials_reducedPartials_sum_40 ^
    reducedPartials_reducedPartials_carry_51 ^ reducedPartials_reducedPartials_carry_50; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_56 = reducedPartials_reducedPartials_sum_40 &
    reducedPartials_reducedPartials_carry_51 | reducedPartials_reducedPartials_carry_51 &
    reducedPartials_reducedPartials_carry_50 | reducedPartials_reducedPartials_sum_40 &
    reducedPartials_reducedPartials_carry_50; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_42 = reducedPartials_reducedPartials_sum_41 ^
    reducedPartials_reducedPartials_carry_49 ^ reducedPartials_reducedPartials_carry_48; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_57 = reducedPartials_reducedPartials_sum_41 &
    reducedPartials_reducedPartials_carry_49 | reducedPartials_reducedPartials_carry_49 &
    reducedPartials_reducedPartials_carry_48 | reducedPartials_reducedPartials_sum_41 &
    reducedPartials_reducedPartials_carry_48; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_43 = reducedPartials_reducedPartials_sum_42 ^
    reducedPartials_reducedPartials_carry_47 ^ partials_27_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_58 = reducedPartials_reducedPartials_sum_42 &
    reducedPartials_reducedPartials_carry_47 | reducedPartials_reducedPartials_carry_47 & partials_27_0 |
    reducedPartials_reducedPartials_sum_42 & partials_27_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_44 = reducedPartials_reducedPartials_sum_43 ^ partials_27_1 ^ partials_27_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_59 = reducedPartials_reducedPartials_sum_43 & partials_27_1 |
    partials_27_1 & partials_27_2 | reducedPartials_reducedPartials_sum_43 & partials_27_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_45 = reducedPartials_reducedPartials_sum_44 ^ partials_27_3 ^ partials_27_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_60 = reducedPartials_reducedPartials_sum_44 & partials_27_3 |
    partials_27_3 & partials_27_4 | reducedPartials_reducedPartials_sum_44 & partials_27_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_46 = reducedPartials_reducedPartials_sum_45 ^ partials_27_5 ^ partials_27_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_61 = reducedPartials_reducedPartials_sum_45 & partials_27_5 |
    partials_27_5 & partials_27_6 | reducedPartials_reducedPartials_sum_45 & partials_27_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_47 = reducedPartials_reducedPartials_sum_46 ^ partials_27_7 ^ partials_27_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_62 = reducedPartials_reducedPartials_sum_46 & partials_27_7 |
    partials_27_7 & partials_27_8 | reducedPartials_reducedPartials_sum_46 & partials_27_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_27_0 = reducedPartials_reducedPartials_sum_47 ^ partials_27_9; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_63 = reducedPartials_reducedPartials_sum_47 & partials_27_9; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_48 = reducedPartials_reducedPartials_carry_63 ^
    reducedPartials_reducedPartials_carry_62 ^ reducedPartials_reducedPartials_carry_61; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_64 = reducedPartials_reducedPartials_carry_63 &
    reducedPartials_reducedPartials_carry_62 | reducedPartials_reducedPartials_carry_62 &
    reducedPartials_reducedPartials_carry_61 | reducedPartials_reducedPartials_carry_63 &
    reducedPartials_reducedPartials_carry_61; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_49 = reducedPartials_reducedPartials_sum_48 ^
    reducedPartials_reducedPartials_carry_60 ^ reducedPartials_reducedPartials_carry_59; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_65 = reducedPartials_reducedPartials_sum_48 &
    reducedPartials_reducedPartials_carry_60 | reducedPartials_reducedPartials_carry_60 &
    reducedPartials_reducedPartials_carry_59 | reducedPartials_reducedPartials_sum_48 &
    reducedPartials_reducedPartials_carry_59; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_50 = reducedPartials_reducedPartials_sum_49 ^
    reducedPartials_reducedPartials_carry_58 ^ reducedPartials_reducedPartials_carry_57; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_66 = reducedPartials_reducedPartials_sum_49 &
    reducedPartials_reducedPartials_carry_58 | reducedPartials_reducedPartials_carry_58 &
    reducedPartials_reducedPartials_carry_57 | reducedPartials_reducedPartials_sum_49 &
    reducedPartials_reducedPartials_carry_57; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_51 = reducedPartials_reducedPartials_sum_50 ^
    reducedPartials_reducedPartials_carry_56 ^ reducedPartials_reducedPartials_carry_55; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_67 = reducedPartials_reducedPartials_sum_50 &
    reducedPartials_reducedPartials_carry_56 | reducedPartials_reducedPartials_carry_56 &
    reducedPartials_reducedPartials_carry_55 | reducedPartials_reducedPartials_sum_50 &
    reducedPartials_reducedPartials_carry_55; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_52 = reducedPartials_reducedPartials_sum_51 ^
    reducedPartials_reducedPartials_28_0 ^ partials_28_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_68 = reducedPartials_reducedPartials_sum_51 &
    reducedPartials_reducedPartials_28_0 | reducedPartials_reducedPartials_28_0 & partials_28_2 |
    reducedPartials_reducedPartials_sum_51 & partials_28_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_53 = reducedPartials_reducedPartials_sum_52 ^ partials_28_3 ^ partials_28_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_69 = reducedPartials_reducedPartials_sum_52 & partials_28_3 |
    partials_28_3 & partials_28_4 | reducedPartials_reducedPartials_sum_52 & partials_28_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_54 = reducedPartials_reducedPartials_sum_53 ^ partials_28_5 ^ partials_28_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_70 = reducedPartials_reducedPartials_sum_53 & partials_28_5 |
    partials_28_5 & partials_28_6 | reducedPartials_reducedPartials_sum_53 & partials_28_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_55 = reducedPartials_reducedPartials_sum_54 ^ partials_28_7 ^ partials_28_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_71 = reducedPartials_reducedPartials_sum_54 & partials_28_7 |
    partials_28_7 & partials_28_8 | reducedPartials_reducedPartials_sum_54 & partials_28_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_28_0_1 = reducedPartials_reducedPartials_sum_55 ^ partials_28_9 ^ partials_28_10
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_72 = reducedPartials_reducedPartials_sum_55 & partials_28_9 |
    partials_28_9 & partials_28_10 | reducedPartials_reducedPartials_sum_55 & partials_28_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_56 = reducedPartials_reducedPartials_carry_72 ^
    reducedPartials_reducedPartials_carry_71 ^ reducedPartials_reducedPartials_carry_70; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_73 = reducedPartials_reducedPartials_carry_72 &
    reducedPartials_reducedPartials_carry_71 | reducedPartials_reducedPartials_carry_71 &
    reducedPartials_reducedPartials_carry_70 | reducedPartials_reducedPartials_carry_72 &
    reducedPartials_reducedPartials_carry_70; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_57 = reducedPartials_reducedPartials_sum_56 ^
    reducedPartials_reducedPartials_carry_69 ^ reducedPartials_reducedPartials_carry_68; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_74 = reducedPartials_reducedPartials_sum_56 &
    reducedPartials_reducedPartials_carry_69 | reducedPartials_reducedPartials_carry_69 &
    reducedPartials_reducedPartials_carry_68 | reducedPartials_reducedPartials_sum_56 &
    reducedPartials_reducedPartials_carry_68; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_58 = reducedPartials_reducedPartials_sum_57 ^
    reducedPartials_reducedPartials_carry_67 ^ reducedPartials_reducedPartials_carry_66; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_75 = reducedPartials_reducedPartials_sum_57 &
    reducedPartials_reducedPartials_carry_67 | reducedPartials_reducedPartials_carry_67 &
    reducedPartials_reducedPartials_carry_66 | reducedPartials_reducedPartials_sum_57 &
    reducedPartials_reducedPartials_carry_66; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_59 = reducedPartials_reducedPartials_sum_58 ^
    reducedPartials_reducedPartials_carry_65 ^ reducedPartials_reducedPartials_carry_64; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_76 = reducedPartials_reducedPartials_sum_58 &
    reducedPartials_reducedPartials_carry_65 | reducedPartials_reducedPartials_carry_65 &
    reducedPartials_reducedPartials_carry_64 | reducedPartials_reducedPartials_sum_58 &
    reducedPartials_reducedPartials_carry_64; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_60 = reducedPartials_reducedPartials_sum_59 ^
    reducedPartials_reducedPartials_29_0 ^ partials_29_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_77 = reducedPartials_reducedPartials_sum_59 &
    reducedPartials_reducedPartials_29_0 | reducedPartials_reducedPartials_29_0 & partials_29_3 |
    reducedPartials_reducedPartials_sum_59 & partials_29_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_61 = reducedPartials_reducedPartials_sum_60 ^ partials_29_4 ^ partials_29_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_78 = reducedPartials_reducedPartials_sum_60 & partials_29_4 |
    partials_29_4 & partials_29_5 | reducedPartials_reducedPartials_sum_60 & partials_29_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_62 = reducedPartials_reducedPartials_sum_61 ^ partials_29_6 ^ partials_29_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_79 = reducedPartials_reducedPartials_sum_61 & partials_29_6 |
    partials_29_6 & partials_29_7 | reducedPartials_reducedPartials_sum_61 & partials_29_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_63 = reducedPartials_reducedPartials_sum_62 ^ partials_29_8 ^ partials_29_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_80 = reducedPartials_reducedPartials_sum_62 & partials_29_8 |
    partials_29_8 & partials_29_9 | reducedPartials_reducedPartials_sum_62 & partials_29_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_29_0_1 = reducedPartials_reducedPartials_sum_63 ^ partials_29_10 ^
    partials_29_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_81 = reducedPartials_reducedPartials_sum_63 & partials_29_10 |
    partials_29_10 & partials_29_11 | reducedPartials_reducedPartials_sum_63 & partials_29_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_64 = reducedPartials_reducedPartials_carry_81 ^
    reducedPartials_reducedPartials_carry_80 ^ reducedPartials_reducedPartials_carry_79; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_82 = reducedPartials_reducedPartials_carry_81 &
    reducedPartials_reducedPartials_carry_80 | reducedPartials_reducedPartials_carry_80 &
    reducedPartials_reducedPartials_carry_79 | reducedPartials_reducedPartials_carry_81 &
    reducedPartials_reducedPartials_carry_79; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_65 = reducedPartials_reducedPartials_sum_64 ^
    reducedPartials_reducedPartials_carry_78 ^ reducedPartials_reducedPartials_carry_77; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_83 = reducedPartials_reducedPartials_sum_64 &
    reducedPartials_reducedPartials_carry_78 | reducedPartials_reducedPartials_carry_78 &
    reducedPartials_reducedPartials_carry_77 | reducedPartials_reducedPartials_sum_64 &
    reducedPartials_reducedPartials_carry_77; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_66 = reducedPartials_reducedPartials_sum_65 ^
    reducedPartials_reducedPartials_carry_76 ^ reducedPartials_reducedPartials_carry_75; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_84 = reducedPartials_reducedPartials_sum_65 &
    reducedPartials_reducedPartials_carry_76 | reducedPartials_reducedPartials_carry_76 &
    reducedPartials_reducedPartials_carry_75 | reducedPartials_reducedPartials_sum_65 &
    reducedPartials_reducedPartials_carry_75; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_67 = reducedPartials_reducedPartials_sum_66 ^
    reducedPartials_reducedPartials_carry_74 ^ reducedPartials_reducedPartials_carry_73; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_85 = reducedPartials_reducedPartials_sum_66 &
    reducedPartials_reducedPartials_carry_74 | reducedPartials_reducedPartials_carry_74 &
    reducedPartials_reducedPartials_carry_73 | reducedPartials_reducedPartials_sum_66 &
    reducedPartials_reducedPartials_carry_73; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_68 = reducedPartials_reducedPartials_sum_67 ^
    reducedPartials_reducedPartials_30_0 ^ partials_30_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_86 = reducedPartials_reducedPartials_sum_67 &
    reducedPartials_reducedPartials_30_0 | reducedPartials_reducedPartials_30_0 & partials_30_4 |
    reducedPartials_reducedPartials_sum_67 & partials_30_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_69 = reducedPartials_reducedPartials_sum_68 ^ partials_30_5 ^ partials_30_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_87 = reducedPartials_reducedPartials_sum_68 & partials_30_5 |
    partials_30_5 & partials_30_6 | reducedPartials_reducedPartials_sum_68 & partials_30_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_70 = reducedPartials_reducedPartials_sum_69 ^ partials_30_7 ^ partials_30_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_88 = reducedPartials_reducedPartials_sum_69 & partials_30_7 |
    partials_30_7 & partials_30_8 | reducedPartials_reducedPartials_sum_69 & partials_30_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_71 = reducedPartials_reducedPartials_sum_70 ^ partials_30_9 ^ partials_30_10
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_89 = reducedPartials_reducedPartials_sum_70 & partials_30_9 |
    partials_30_9 & partials_30_10 | reducedPartials_reducedPartials_sum_70 & partials_30_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_30_0_1 = reducedPartials_reducedPartials_sum_71 ^ partials_30_11 ^
    partials_30_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_90 = reducedPartials_reducedPartials_sum_71 & partials_30_11 |
    partials_30_11 & partials_30_12 | reducedPartials_reducedPartials_sum_71 & partials_30_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_72 = reducedPartials_reducedPartials_carry_90 ^
    reducedPartials_reducedPartials_carry_89 ^ reducedPartials_reducedPartials_carry_88; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_91 = reducedPartials_reducedPartials_carry_90 &
    reducedPartials_reducedPartials_carry_89 | reducedPartials_reducedPartials_carry_89 &
    reducedPartials_reducedPartials_carry_88 | reducedPartials_reducedPartials_carry_90 &
    reducedPartials_reducedPartials_carry_88; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_73 = reducedPartials_reducedPartials_sum_72 ^
    reducedPartials_reducedPartials_carry_87 ^ reducedPartials_reducedPartials_carry_86; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_92 = reducedPartials_reducedPartials_sum_72 &
    reducedPartials_reducedPartials_carry_87 | reducedPartials_reducedPartials_carry_87 &
    reducedPartials_reducedPartials_carry_86 | reducedPartials_reducedPartials_sum_72 &
    reducedPartials_reducedPartials_carry_86; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_74 = reducedPartials_reducedPartials_sum_73 ^
    reducedPartials_reducedPartials_carry_85 ^ reducedPartials_reducedPartials_carry_84; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_93 = reducedPartials_reducedPartials_sum_73 &
    reducedPartials_reducedPartials_carry_85 | reducedPartials_reducedPartials_carry_85 &
    reducedPartials_reducedPartials_carry_84 | reducedPartials_reducedPartials_sum_73 &
    reducedPartials_reducedPartials_carry_84; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_75 = reducedPartials_reducedPartials_sum_74 ^
    reducedPartials_reducedPartials_carry_83 ^ reducedPartials_reducedPartials_carry_82; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_94 = reducedPartials_reducedPartials_sum_74 &
    reducedPartials_reducedPartials_carry_83 | reducedPartials_reducedPartials_carry_83 &
    reducedPartials_reducedPartials_carry_82 | reducedPartials_reducedPartials_sum_74 &
    reducedPartials_reducedPartials_carry_82; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_76 = reducedPartials_reducedPartials_sum_75 ^
    reducedPartials_reducedPartials_31_0 ^ partials_31_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_95 = reducedPartials_reducedPartials_sum_75 &
    reducedPartials_reducedPartials_31_0 | reducedPartials_reducedPartials_31_0 & partials_31_5 |
    reducedPartials_reducedPartials_sum_75 & partials_31_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_77 = reducedPartials_reducedPartials_sum_76 ^ partials_31_6 ^ partials_31_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_96 = reducedPartials_reducedPartials_sum_76 & partials_31_6 |
    partials_31_6 & partials_31_7 | reducedPartials_reducedPartials_sum_76 & partials_31_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_78 = reducedPartials_reducedPartials_sum_77 ^ partials_31_8 ^ partials_31_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_97 = reducedPartials_reducedPartials_sum_77 & partials_31_8 |
    partials_31_8 & partials_31_9 | reducedPartials_reducedPartials_sum_77 & partials_31_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_79 = reducedPartials_reducedPartials_sum_78 ^ partials_31_10 ^
    partials_31_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_98 = reducedPartials_reducedPartials_sum_78 & partials_31_10 |
    partials_31_10 & partials_31_11 | reducedPartials_reducedPartials_sum_78 & partials_31_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_31_0_1 = reducedPartials_reducedPartials_sum_79 ^ partials_31_12 ^
    partials_31_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_99 = reducedPartials_reducedPartials_sum_79 & partials_31_12 |
    partials_31_12 & partials_31_13 | reducedPartials_reducedPartials_sum_79 & partials_31_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_80 = reducedPartials_reducedPartials_carry_99 ^
    reducedPartials_reducedPartials_carry_98 ^ reducedPartials_reducedPartials_carry_97; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_100 = reducedPartials_reducedPartials_carry_99 &
    reducedPartials_reducedPartials_carry_98 | reducedPartials_reducedPartials_carry_98 &
    reducedPartials_reducedPartials_carry_97 | reducedPartials_reducedPartials_carry_99 &
    reducedPartials_reducedPartials_carry_97; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_81 = reducedPartials_reducedPartials_sum_80 ^
    reducedPartials_reducedPartials_carry_96 ^ reducedPartials_reducedPartials_carry_95; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_101 = reducedPartials_reducedPartials_sum_80 &
    reducedPartials_reducedPartials_carry_96 | reducedPartials_reducedPartials_carry_96 &
    reducedPartials_reducedPartials_carry_95 | reducedPartials_reducedPartials_sum_80 &
    reducedPartials_reducedPartials_carry_95; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_82 = reducedPartials_reducedPartials_sum_81 ^
    reducedPartials_reducedPartials_carry_94 ^ reducedPartials_reducedPartials_carry_93; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_102 = reducedPartials_reducedPartials_sum_81 &
    reducedPartials_reducedPartials_carry_94 | reducedPartials_reducedPartials_carry_94 &
    reducedPartials_reducedPartials_carry_93 | reducedPartials_reducedPartials_sum_81 &
    reducedPartials_reducedPartials_carry_93; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_83 = reducedPartials_reducedPartials_sum_82 ^
    reducedPartials_reducedPartials_carry_92 ^ reducedPartials_reducedPartials_carry_91; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_103 = reducedPartials_reducedPartials_sum_82 &
    reducedPartials_reducedPartials_carry_92 | reducedPartials_reducedPartials_carry_92 &
    reducedPartials_reducedPartials_carry_91 | reducedPartials_reducedPartials_sum_82 &
    reducedPartials_reducedPartials_carry_91; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_84 = reducedPartials_reducedPartials_sum_83 ^
    reducedPartials_reducedPartials_32_0 ^ partials_32_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_104 = reducedPartials_reducedPartials_sum_83 &
    reducedPartials_reducedPartials_32_0 | reducedPartials_reducedPartials_32_0 & partials_32_4 |
    reducedPartials_reducedPartials_sum_83 & partials_32_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_85 = reducedPartials_reducedPartials_sum_84 ^ partials_32_5 ^ partials_32_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_105 = reducedPartials_reducedPartials_sum_84 & partials_32_5 |
    partials_32_5 & partials_32_6 | reducedPartials_reducedPartials_sum_84 & partials_32_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_86 = reducedPartials_reducedPartials_sum_85 ^ partials_32_7 ^ partials_32_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_106 = reducedPartials_reducedPartials_sum_85 & partials_32_7 |
    partials_32_7 & partials_32_8 | reducedPartials_reducedPartials_sum_85 & partials_32_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_87 = reducedPartials_reducedPartials_sum_86 ^ partials_32_9 ^ partials_32_10
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_107 = reducedPartials_reducedPartials_sum_86 & partials_32_9 |
    partials_32_9 & partials_32_10 | reducedPartials_reducedPartials_sum_86 & partials_32_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_32_0_1 = reducedPartials_reducedPartials_sum_87 ^ partials_32_11 ^
    partials_32_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_108 = reducedPartials_reducedPartials_sum_87 & partials_32_11 |
    partials_32_11 & partials_32_12 | reducedPartials_reducedPartials_sum_87 & partials_32_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_88 = reducedPartials_reducedPartials_carry_108 ^
    reducedPartials_reducedPartials_carry_107 ^ reducedPartials_reducedPartials_carry_106; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_109 = reducedPartials_reducedPartials_carry_108 &
    reducedPartials_reducedPartials_carry_107 | reducedPartials_reducedPartials_carry_107 &
    reducedPartials_reducedPartials_carry_106 | reducedPartials_reducedPartials_carry_108 &
    reducedPartials_reducedPartials_carry_106; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_89 = reducedPartials_reducedPartials_sum_88 ^
    reducedPartials_reducedPartials_carry_105 ^ reducedPartials_reducedPartials_carry_104; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_110 = reducedPartials_reducedPartials_sum_88 &
    reducedPartials_reducedPartials_carry_105 | reducedPartials_reducedPartials_carry_105 &
    reducedPartials_reducedPartials_carry_104 | reducedPartials_reducedPartials_sum_88 &
    reducedPartials_reducedPartials_carry_104; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_90 = reducedPartials_reducedPartials_sum_89 ^
    reducedPartials_reducedPartials_carry_103 ^ reducedPartials_reducedPartials_carry_102; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_111 = reducedPartials_reducedPartials_sum_89 &
    reducedPartials_reducedPartials_carry_103 | reducedPartials_reducedPartials_carry_103 &
    reducedPartials_reducedPartials_carry_102 | reducedPartials_reducedPartials_sum_89 &
    reducedPartials_reducedPartials_carry_102; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_91 = reducedPartials_reducedPartials_sum_90 ^
    reducedPartials_reducedPartials_carry_101 ^ reducedPartials_reducedPartials_carry_100; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_112 = reducedPartials_reducedPartials_sum_90 &
    reducedPartials_reducedPartials_carry_101 | reducedPartials_reducedPartials_carry_101 &
    reducedPartials_reducedPartials_carry_100 | reducedPartials_reducedPartials_sum_90 &
    reducedPartials_reducedPartials_carry_100; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_92 = reducedPartials_reducedPartials_sum_91 ^
    reducedPartials_reducedPartials_33_0 ^ partials_33_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_113 = reducedPartials_reducedPartials_sum_91 &
    reducedPartials_reducedPartials_33_0 | reducedPartials_reducedPartials_33_0 & partials_33_3 |
    reducedPartials_reducedPartials_sum_91 & partials_33_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_93 = reducedPartials_reducedPartials_sum_92 ^ partials_33_4 ^ partials_33_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_114 = reducedPartials_reducedPartials_sum_92 & partials_33_4 |
    partials_33_4 & partials_33_5 | reducedPartials_reducedPartials_sum_92 & partials_33_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_94 = reducedPartials_reducedPartials_sum_93 ^ partials_33_6 ^ partials_33_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_115 = reducedPartials_reducedPartials_sum_93 & partials_33_6 |
    partials_33_6 & partials_33_7 | reducedPartials_reducedPartials_sum_93 & partials_33_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_95 = reducedPartials_reducedPartials_sum_94 ^ partials_33_8 ^ partials_33_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_116 = reducedPartials_reducedPartials_sum_94 & partials_33_8 |
    partials_33_8 & partials_33_9 | reducedPartials_reducedPartials_sum_94 & partials_33_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_33_0_1 = reducedPartials_reducedPartials_sum_95 ^ partials_33_10 ^
    partials_33_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_117 = reducedPartials_reducedPartials_sum_95 & partials_33_10 |
    partials_33_10 & partials_33_11 | reducedPartials_reducedPartials_sum_95 & partials_33_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_96 = reducedPartials_reducedPartials_carry_117 ^
    reducedPartials_reducedPartials_carry_116 ^ reducedPartials_reducedPartials_carry_115; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_118 = reducedPartials_reducedPartials_carry_117 &
    reducedPartials_reducedPartials_carry_116 | reducedPartials_reducedPartials_carry_116 &
    reducedPartials_reducedPartials_carry_115 | reducedPartials_reducedPartials_carry_117 &
    reducedPartials_reducedPartials_carry_115; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_97 = reducedPartials_reducedPartials_sum_96 ^
    reducedPartials_reducedPartials_carry_114 ^ reducedPartials_reducedPartials_carry_113; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_119 = reducedPartials_reducedPartials_sum_96 &
    reducedPartials_reducedPartials_carry_114 | reducedPartials_reducedPartials_carry_114 &
    reducedPartials_reducedPartials_carry_113 | reducedPartials_reducedPartials_sum_96 &
    reducedPartials_reducedPartials_carry_113; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_98 = reducedPartials_reducedPartials_sum_97 ^
    reducedPartials_reducedPartials_carry_112 ^ reducedPartials_reducedPartials_carry_111; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_120 = reducedPartials_reducedPartials_sum_97 &
    reducedPartials_reducedPartials_carry_112 | reducedPartials_reducedPartials_carry_112 &
    reducedPartials_reducedPartials_carry_111 | reducedPartials_reducedPartials_sum_97 &
    reducedPartials_reducedPartials_carry_111; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_99 = reducedPartials_reducedPartials_sum_98 ^
    reducedPartials_reducedPartials_carry_110 ^ reducedPartials_reducedPartials_carry_109; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_121 = reducedPartials_reducedPartials_sum_98 &
    reducedPartials_reducedPartials_carry_110 | reducedPartials_reducedPartials_carry_110 &
    reducedPartials_reducedPartials_carry_109 | reducedPartials_reducedPartials_sum_98 &
    reducedPartials_reducedPartials_carry_109; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_100 = reducedPartials_reducedPartials_sum_99 ^
    reducedPartials_reducedPartials_34_0 ^ partials_34_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_122 = reducedPartials_reducedPartials_sum_99 &
    reducedPartials_reducedPartials_34_0 | reducedPartials_reducedPartials_34_0 & partials_34_2 |
    reducedPartials_reducedPartials_sum_99 & partials_34_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_101 = reducedPartials_reducedPartials_sum_100 ^ partials_34_3 ^
    partials_34_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_123 = reducedPartials_reducedPartials_sum_100 & partials_34_3 |
    partials_34_3 & partials_34_4 | reducedPartials_reducedPartials_sum_100 & partials_34_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_102 = reducedPartials_reducedPartials_sum_101 ^ partials_34_5 ^
    partials_34_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_124 = reducedPartials_reducedPartials_sum_101 & partials_34_5 |
    partials_34_5 & partials_34_6 | reducedPartials_reducedPartials_sum_101 & partials_34_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_103 = reducedPartials_reducedPartials_sum_102 ^ partials_34_7 ^
    partials_34_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_125 = reducedPartials_reducedPartials_sum_102 & partials_34_7 |
    partials_34_7 & partials_34_8 | reducedPartials_reducedPartials_sum_102 & partials_34_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_34_0_1 = reducedPartials_reducedPartials_sum_103 ^ partials_34_9 ^
    partials_34_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_126 = reducedPartials_reducedPartials_sum_103 & partials_34_9 |
    partials_34_9 & partials_34_10 | reducedPartials_reducedPartials_sum_103 & partials_34_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_104 = reducedPartials_reducedPartials_carry_126 ^
    reducedPartials_reducedPartials_carry_125 ^ reducedPartials_reducedPartials_carry_124; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_127 = reducedPartials_reducedPartials_carry_126 &
    reducedPartials_reducedPartials_carry_125 | reducedPartials_reducedPartials_carry_125 &
    reducedPartials_reducedPartials_carry_124 | reducedPartials_reducedPartials_carry_126 &
    reducedPartials_reducedPartials_carry_124; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_105 = reducedPartials_reducedPartials_sum_104 ^
    reducedPartials_reducedPartials_carry_123 ^ reducedPartials_reducedPartials_carry_122; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_128 = reducedPartials_reducedPartials_sum_104 &
    reducedPartials_reducedPartials_carry_123 | reducedPartials_reducedPartials_carry_123 &
    reducedPartials_reducedPartials_carry_122 | reducedPartials_reducedPartials_sum_104 &
    reducedPartials_reducedPartials_carry_122; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_106 = reducedPartials_reducedPartials_sum_105 ^
    reducedPartials_reducedPartials_carry_121 ^ reducedPartials_reducedPartials_carry_120; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_129 = reducedPartials_reducedPartials_sum_105 &
    reducedPartials_reducedPartials_carry_121 | reducedPartials_reducedPartials_carry_121 &
    reducedPartials_reducedPartials_carry_120 | reducedPartials_reducedPartials_sum_105 &
    reducedPartials_reducedPartials_carry_120; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_107 = reducedPartials_reducedPartials_sum_106 ^
    reducedPartials_reducedPartials_carry_119 ^ reducedPartials_reducedPartials_carry_118; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_130 = reducedPartials_reducedPartials_sum_106 &
    reducedPartials_reducedPartials_carry_119 | reducedPartials_reducedPartials_carry_119 &
    reducedPartials_reducedPartials_carry_118 | reducedPartials_reducedPartials_sum_106 &
    reducedPartials_reducedPartials_carry_118; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_108 = reducedPartials_reducedPartials_sum_107 ^
    reducedPartials_reducedPartials_35_0 ^ partials_35_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_131 = reducedPartials_reducedPartials_sum_107 &
    reducedPartials_reducedPartials_35_0 | reducedPartials_reducedPartials_35_0 & partials_35_1 |
    reducedPartials_reducedPartials_sum_107 & partials_35_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_109 = reducedPartials_reducedPartials_sum_108 ^ partials_35_2 ^
    partials_35_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_132 = reducedPartials_reducedPartials_sum_108 & partials_35_2 |
    partials_35_2 & partials_35_3 | reducedPartials_reducedPartials_sum_108 & partials_35_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_110 = reducedPartials_reducedPartials_sum_109 ^ partials_35_4 ^
    partials_35_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_133 = reducedPartials_reducedPartials_sum_109 & partials_35_4 |
    partials_35_4 & partials_35_5 | reducedPartials_reducedPartials_sum_109 & partials_35_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_111 = reducedPartials_reducedPartials_sum_110 ^ partials_35_6 ^
    partials_35_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_134 = reducedPartials_reducedPartials_sum_110 & partials_35_6 |
    partials_35_6 & partials_35_7 | reducedPartials_reducedPartials_sum_110 & partials_35_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_35_0_1 = reducedPartials_reducedPartials_sum_111 ^ partials_35_8 ^ partials_35_9
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_135 = reducedPartials_reducedPartials_sum_111 & partials_35_8 |
    partials_35_8 & partials_35_9 | reducedPartials_reducedPartials_sum_111 & partials_35_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_112 = reducedPartials_reducedPartials_carry_135 ^
    reducedPartials_reducedPartials_carry_134 ^ reducedPartials_reducedPartials_carry_133; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_136 = reducedPartials_reducedPartials_carry_135 &
    reducedPartials_reducedPartials_carry_134 | reducedPartials_reducedPartials_carry_134 &
    reducedPartials_reducedPartials_carry_133 | reducedPartials_reducedPartials_carry_135 &
    reducedPartials_reducedPartials_carry_133; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_113 = reducedPartials_reducedPartials_sum_112 ^
    reducedPartials_reducedPartials_carry_132 ^ reducedPartials_reducedPartials_carry_131; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_137 = reducedPartials_reducedPartials_sum_112 &
    reducedPartials_reducedPartials_carry_132 | reducedPartials_reducedPartials_carry_132 &
    reducedPartials_reducedPartials_carry_131 | reducedPartials_reducedPartials_sum_112 &
    reducedPartials_reducedPartials_carry_131; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_114 = reducedPartials_reducedPartials_sum_113 ^
    reducedPartials_reducedPartials_carry_130 ^ reducedPartials_reducedPartials_carry_129; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_138 = reducedPartials_reducedPartials_sum_113 &
    reducedPartials_reducedPartials_carry_130 | reducedPartials_reducedPartials_carry_130 &
    reducedPartials_reducedPartials_carry_129 | reducedPartials_reducedPartials_sum_113 &
    reducedPartials_reducedPartials_carry_129; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_115 = reducedPartials_reducedPartials_sum_114 ^
    reducedPartials_reducedPartials_carry_128 ^ reducedPartials_reducedPartials_carry_127; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_139 = reducedPartials_reducedPartials_sum_114 &
    reducedPartials_reducedPartials_carry_128 | reducedPartials_reducedPartials_carry_128 &
    reducedPartials_reducedPartials_carry_127 | reducedPartials_reducedPartials_sum_114 &
    reducedPartials_reducedPartials_carry_127; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_116 = reducedPartials_reducedPartials_sum_115 ^
    reducedPartials_reducedPartials_36_0 ^ partials_36_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_140 = reducedPartials_reducedPartials_sum_115 &
    reducedPartials_reducedPartials_36_0 | reducedPartials_reducedPartials_36_0 & partials_36_0 |
    reducedPartials_reducedPartials_sum_115 & partials_36_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_117 = reducedPartials_reducedPartials_sum_116 ^ partials_36_1 ^
    partials_36_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_141 = reducedPartials_reducedPartials_sum_116 & partials_36_1 |
    partials_36_1 & partials_36_2 | reducedPartials_reducedPartials_sum_116 & partials_36_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_118 = reducedPartials_reducedPartials_sum_117 ^ partials_36_3 ^
    partials_36_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_142 = reducedPartials_reducedPartials_sum_117 & partials_36_3 |
    partials_36_3 & partials_36_4 | reducedPartials_reducedPartials_sum_117 & partials_36_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_119 = reducedPartials_reducedPartials_sum_118 ^ partials_36_5 ^
    partials_36_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_143 = reducedPartials_reducedPartials_sum_118 & partials_36_5 |
    partials_36_5 & partials_36_6 | reducedPartials_reducedPartials_sum_118 & partials_36_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_36_0_1 = reducedPartials_reducedPartials_sum_119 ^ partials_36_7 ^ partials_36_8
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_144 = reducedPartials_reducedPartials_sum_119 & partials_36_7 |
    partials_36_7 & partials_36_8 | reducedPartials_reducedPartials_sum_119 & partials_36_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_120 = reducedPartials_reducedPartials_carry_144 ^
    reducedPartials_reducedPartials_carry_143 ^ reducedPartials_reducedPartials_carry_142; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_145 = reducedPartials_reducedPartials_carry_144 &
    reducedPartials_reducedPartials_carry_143 | reducedPartials_reducedPartials_carry_143 &
    reducedPartials_reducedPartials_carry_142 | reducedPartials_reducedPartials_carry_144 &
    reducedPartials_reducedPartials_carry_142; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_121 = reducedPartials_reducedPartials_sum_120 ^
    reducedPartials_reducedPartials_carry_141 ^ reducedPartials_reducedPartials_carry_140; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_146 = reducedPartials_reducedPartials_sum_120 &
    reducedPartials_reducedPartials_carry_141 | reducedPartials_reducedPartials_carry_141 &
    reducedPartials_reducedPartials_carry_140 | reducedPartials_reducedPartials_sum_120 &
    reducedPartials_reducedPartials_carry_140; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_122 = reducedPartials_reducedPartials_sum_121 ^
    reducedPartials_reducedPartials_carry_139 ^ reducedPartials_reducedPartials_carry_138; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_147 = reducedPartials_reducedPartials_sum_121 &
    reducedPartials_reducedPartials_carry_139 | reducedPartials_reducedPartials_carry_139 &
    reducedPartials_reducedPartials_carry_138 | reducedPartials_reducedPartials_sum_121 &
    reducedPartials_reducedPartials_carry_138; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_123 = reducedPartials_reducedPartials_sum_122 ^
    reducedPartials_reducedPartials_carry_137 ^ reducedPartials_reducedPartials_carry_136; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_148 = reducedPartials_reducedPartials_sum_122 &
    reducedPartials_reducedPartials_carry_137 | reducedPartials_reducedPartials_carry_137 &
    reducedPartials_reducedPartials_carry_136 | reducedPartials_reducedPartials_sum_122 &
    reducedPartials_reducedPartials_carry_136; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_124 = reducedPartials_reducedPartials_sum_123 ^ partials_37_0 ^
    partials_37_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_149 = reducedPartials_reducedPartials_sum_123 & partials_37_0 |
    partials_37_0 & partials_37_1 | reducedPartials_reducedPartials_sum_123 & partials_37_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_125 = reducedPartials_reducedPartials_sum_124 ^ partials_37_2 ^
    partials_37_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_150 = reducedPartials_reducedPartials_sum_124 & partials_37_2 |
    partials_37_2 & partials_37_3 | reducedPartials_reducedPartials_sum_124 & partials_37_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_126 = reducedPartials_reducedPartials_sum_125 ^ partials_37_4 ^
    partials_37_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_151 = reducedPartials_reducedPartials_sum_125 & partials_37_4 |
    partials_37_4 & partials_37_5 | reducedPartials_reducedPartials_sum_125 & partials_37_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_37_0 = reducedPartials_reducedPartials_sum_126 ^ partials_37_6 ^ partials_37_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_152 = reducedPartials_reducedPartials_sum_126 & partials_37_6 |
    partials_37_6 & partials_37_7 | reducedPartials_reducedPartials_sum_126 & partials_37_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_127 = reducedPartials_reducedPartials_carry_152 ^
    reducedPartials_reducedPartials_carry_151 ^ reducedPartials_reducedPartials_carry_150; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_153 = reducedPartials_reducedPartials_carry_152 &
    reducedPartials_reducedPartials_carry_151 | reducedPartials_reducedPartials_carry_151 &
    reducedPartials_reducedPartials_carry_150 | reducedPartials_reducedPartials_carry_152 &
    reducedPartials_reducedPartials_carry_150; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_128 = reducedPartials_reducedPartials_sum_127 ^
    reducedPartials_reducedPartials_carry_149 ^ reducedPartials_reducedPartials_carry_148; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_154 = reducedPartials_reducedPartials_sum_127 &
    reducedPartials_reducedPartials_carry_149 | reducedPartials_reducedPartials_carry_149 &
    reducedPartials_reducedPartials_carry_148 | reducedPartials_reducedPartials_sum_127 &
    reducedPartials_reducedPartials_carry_148; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_129 = reducedPartials_reducedPartials_sum_128 ^
    reducedPartials_reducedPartials_carry_147 ^ reducedPartials_reducedPartials_carry_146; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_155 = reducedPartials_reducedPartials_sum_128 &
    reducedPartials_reducedPartials_carry_147 | reducedPartials_reducedPartials_carry_147 &
    reducedPartials_reducedPartials_carry_146 | reducedPartials_reducedPartials_sum_128 &
    reducedPartials_reducedPartials_carry_146; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_130 = reducedPartials_reducedPartials_sum_129 ^
    reducedPartials_reducedPartials_carry_145 ^ partials_38_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_156 = reducedPartials_reducedPartials_sum_129 &
    reducedPartials_reducedPartials_carry_145 | reducedPartials_reducedPartials_carry_145 & partials_38_0 |
    reducedPartials_reducedPartials_sum_129 & partials_38_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_131 = reducedPartials_reducedPartials_sum_130 ^ partials_38_1 ^
    partials_38_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_157 = reducedPartials_reducedPartials_sum_130 & partials_38_1 |
    partials_38_1 & partials_38_2 | reducedPartials_reducedPartials_sum_130 & partials_38_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_132 = reducedPartials_reducedPartials_sum_131 ^ partials_38_3 ^
    partials_38_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_158 = reducedPartials_reducedPartials_sum_131 & partials_38_3 |
    partials_38_3 & partials_38_4 | reducedPartials_reducedPartials_sum_131 & partials_38_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_38_0 = reducedPartials_reducedPartials_sum_132 ^ partials_38_5 ^ partials_38_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_159 = reducedPartials_reducedPartials_sum_132 & partials_38_5 |
    partials_38_5 & partials_38_6 | reducedPartials_reducedPartials_sum_132 & partials_38_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_133 = reducedPartials_reducedPartials_carry_159 ^
    reducedPartials_reducedPartials_carry_158 ^ reducedPartials_reducedPartials_carry_157; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_160 = reducedPartials_reducedPartials_carry_159 &
    reducedPartials_reducedPartials_carry_158 | reducedPartials_reducedPartials_carry_158 &
    reducedPartials_reducedPartials_carry_157 | reducedPartials_reducedPartials_carry_159 &
    reducedPartials_reducedPartials_carry_157; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_134 = reducedPartials_reducedPartials_sum_133 ^
    reducedPartials_reducedPartials_carry_156 ^ reducedPartials_reducedPartials_carry_155; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_161 = reducedPartials_reducedPartials_sum_133 &
    reducedPartials_reducedPartials_carry_156 | reducedPartials_reducedPartials_carry_156 &
    reducedPartials_reducedPartials_carry_155 | reducedPartials_reducedPartials_sum_133 &
    reducedPartials_reducedPartials_carry_155; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_135 = reducedPartials_reducedPartials_sum_134 ^
    reducedPartials_reducedPartials_carry_154 ^ reducedPartials_reducedPartials_carry_153; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_162 = reducedPartials_reducedPartials_sum_134 &
    reducedPartials_reducedPartials_carry_154 | reducedPartials_reducedPartials_carry_154 &
    reducedPartials_reducedPartials_carry_153 | reducedPartials_reducedPartials_sum_134 &
    reducedPartials_reducedPartials_carry_153; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_136 = reducedPartials_reducedPartials_sum_135 ^ partials_39_0 ^
    partials_39_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_163 = reducedPartials_reducedPartials_sum_135 & partials_39_0 |
    partials_39_0 & partials_39_1 | reducedPartials_reducedPartials_sum_135 & partials_39_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_137 = reducedPartials_reducedPartials_sum_136 ^ partials_39_2 ^
    partials_39_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_164 = reducedPartials_reducedPartials_sum_136 & partials_39_2 |
    partials_39_2 & partials_39_3 | reducedPartials_reducedPartials_sum_136 & partials_39_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_39_0 = reducedPartials_reducedPartials_sum_137 ^ partials_39_4 ^ partials_39_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_165 = reducedPartials_reducedPartials_sum_137 & partials_39_4 |
    partials_39_4 & partials_39_5 | reducedPartials_reducedPartials_sum_137 & partials_39_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_138 = reducedPartials_reducedPartials_carry_165 ^
    reducedPartials_reducedPartials_carry_164 ^ reducedPartials_reducedPartials_carry_163; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_166 = reducedPartials_reducedPartials_carry_165 &
    reducedPartials_reducedPartials_carry_164 | reducedPartials_reducedPartials_carry_164 &
    reducedPartials_reducedPartials_carry_163 | reducedPartials_reducedPartials_carry_165 &
    reducedPartials_reducedPartials_carry_163; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_139 = reducedPartials_reducedPartials_sum_138 ^
    reducedPartials_reducedPartials_carry_162 ^ reducedPartials_reducedPartials_carry_161; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_167 = reducedPartials_reducedPartials_sum_138 &
    reducedPartials_reducedPartials_carry_162 | reducedPartials_reducedPartials_carry_162 &
    reducedPartials_reducedPartials_carry_161 | reducedPartials_reducedPartials_sum_138 &
    reducedPartials_reducedPartials_carry_161; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_140 = reducedPartials_reducedPartials_sum_139 ^
    reducedPartials_reducedPartials_carry_160 ^ partials_40_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_168 = reducedPartials_reducedPartials_sum_139 &
    reducedPartials_reducedPartials_carry_160 | reducedPartials_reducedPartials_carry_160 & partials_40_0 |
    reducedPartials_reducedPartials_sum_139 & partials_40_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_141 = reducedPartials_reducedPartials_sum_140 ^ partials_40_1 ^
    partials_40_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_169 = reducedPartials_reducedPartials_sum_140 & partials_40_1 |
    partials_40_1 & partials_40_2 | reducedPartials_reducedPartials_sum_140 & partials_40_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_40_0 = reducedPartials_reducedPartials_sum_141 ^ partials_40_3 ^ partials_40_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_170 = reducedPartials_reducedPartials_sum_141 & partials_40_3 |
    partials_40_3 & partials_40_4 | reducedPartials_reducedPartials_sum_141 & partials_40_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_142 = reducedPartials_reducedPartials_carry_170 ^
    reducedPartials_reducedPartials_carry_169 ^ reducedPartials_reducedPartials_carry_168; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_171 = reducedPartials_reducedPartials_carry_170 &
    reducedPartials_reducedPartials_carry_169 | reducedPartials_reducedPartials_carry_169 &
    reducedPartials_reducedPartials_carry_168 | reducedPartials_reducedPartials_carry_170 &
    reducedPartials_reducedPartials_carry_168; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_143 = reducedPartials_reducedPartials_sum_142 ^
    reducedPartials_reducedPartials_carry_167 ^ reducedPartials_reducedPartials_carry_166; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_172 = reducedPartials_reducedPartials_sum_142 &
    reducedPartials_reducedPartials_carry_167 | reducedPartials_reducedPartials_carry_167 &
    reducedPartials_reducedPartials_carry_166 | reducedPartials_reducedPartials_sum_142 &
    reducedPartials_reducedPartials_carry_166; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_144 = reducedPartials_reducedPartials_sum_143 ^ partials_41_0 ^
    partials_41_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_173 = reducedPartials_reducedPartials_sum_143 & partials_41_0 |
    partials_41_0 & partials_41_1 | reducedPartials_reducedPartials_sum_143 & partials_41_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_41_0 = reducedPartials_reducedPartials_sum_144 ^ partials_41_2 ^ partials_41_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_174 = reducedPartials_reducedPartials_sum_144 & partials_41_2 |
    partials_41_2 & partials_41_3 | reducedPartials_reducedPartials_sum_144 & partials_41_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_145 = reducedPartials_reducedPartials_carry_174 ^
    reducedPartials_reducedPartials_carry_173 ^ reducedPartials_reducedPartials_carry_172; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_175 = reducedPartials_reducedPartials_carry_174 &
    reducedPartials_reducedPartials_carry_173 | reducedPartials_reducedPartials_carry_173 &
    reducedPartials_reducedPartials_carry_172 | reducedPartials_reducedPartials_carry_174 &
    reducedPartials_reducedPartials_carry_172; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_146 = reducedPartials_reducedPartials_sum_145 ^
    reducedPartials_reducedPartials_carry_171 ^ partials_42_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_176 = reducedPartials_reducedPartials_sum_145 &
    reducedPartials_reducedPartials_carry_171 | reducedPartials_reducedPartials_carry_171 & partials_42_0 |
    reducedPartials_reducedPartials_sum_145 & partials_42_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_42_0 = reducedPartials_reducedPartials_sum_146 ^ partials_42_1 ^ partials_42_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_177 = reducedPartials_reducedPartials_sum_146 & partials_42_1 |
    partials_42_1 & partials_42_2 | reducedPartials_reducedPartials_sum_146 & partials_42_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_147 = reducedPartials_reducedPartials_carry_177 ^
    reducedPartials_reducedPartials_carry_176 ^ reducedPartials_reducedPartials_carry_175; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_178 = reducedPartials_reducedPartials_carry_177 &
    reducedPartials_reducedPartials_carry_176 | reducedPartials_reducedPartials_carry_176 &
    reducedPartials_reducedPartials_carry_175 | reducedPartials_reducedPartials_carry_177 &
    reducedPartials_reducedPartials_carry_175; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_43_0 = reducedPartials_reducedPartials_sum_147 ^ partials_43_0 ^ partials_43_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_179 = reducedPartials_reducedPartials_sum_147 & partials_43_0 |
    partials_43_0 & partials_43_1 | reducedPartials_reducedPartials_sum_147 & partials_43_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_44_0 = reducedPartials_reducedPartials_carry_179 ^
    reducedPartials_reducedPartials_carry_178 ^ partials_44_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_45_0 = reducedPartials_reducedPartials_carry_179 &
    reducedPartials_reducedPartials_carry_178 | reducedPartials_reducedPartials_carry_178 & partials_44_0 |
    reducedPartials_reducedPartials_carry_179 & partials_44_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_13_0 = partials_13_0 ^ partials_13_1; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_180 = partials_13_0 & partials_13_1; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_148 = reducedPartials_reducedPartials_carry_180 ^ partials_14_0 ^
    partials_14_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_181 = reducedPartials_reducedPartials_carry_180 & partials_14_0 |
    partials_14_0 & partials_14_1 | reducedPartials_reducedPartials_carry_180 & partials_14_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_14_0 = reducedPartials_reducedPartials_sum_148 ^ partials_14_2; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_182 = reducedPartials_reducedPartials_sum_148 & partials_14_2; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_149 = reducedPartials_reducedPartials_carry_182 ^
    reducedPartials_reducedPartials_carry_181 ^ partials_15_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_183 = reducedPartials_reducedPartials_carry_182 &
    reducedPartials_reducedPartials_carry_181 | reducedPartials_reducedPartials_carry_181 & partials_15_0 |
    reducedPartials_reducedPartials_carry_182 & partials_15_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_150 = reducedPartials_reducedPartials_sum_149 ^ partials_15_1 ^
    partials_15_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_184 = reducedPartials_reducedPartials_sum_149 & partials_15_1 |
    partials_15_1 & partials_15_2 | reducedPartials_reducedPartials_sum_149 & partials_15_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_15_0 = reducedPartials_reducedPartials_sum_150 ^ partials_15_3; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_185 = reducedPartials_reducedPartials_sum_150 & partials_15_3; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_151 = reducedPartials_reducedPartials_carry_185 ^
    reducedPartials_reducedPartials_carry_184 ^ reducedPartials_reducedPartials_carry_183; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_186 = reducedPartials_reducedPartials_carry_185 &
    reducedPartials_reducedPartials_carry_184 | reducedPartials_reducedPartials_carry_184 &
    reducedPartials_reducedPartials_carry_183 | reducedPartials_reducedPartials_carry_185 &
    reducedPartials_reducedPartials_carry_183; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_152 = reducedPartials_reducedPartials_sum_151 ^ partials_16_0 ^
    partials_16_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_187 = reducedPartials_reducedPartials_sum_151 & partials_16_0 |
    partials_16_0 & partials_16_1 | reducedPartials_reducedPartials_sum_151 & partials_16_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_153 = reducedPartials_reducedPartials_sum_152 ^ partials_16_2 ^
    partials_16_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_188 = reducedPartials_reducedPartials_sum_152 & partials_16_2 |
    partials_16_2 & partials_16_3 | reducedPartials_reducedPartials_sum_152 & partials_16_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_16_0 = reducedPartials_reducedPartials_sum_153 ^ partials_16_4; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_189 = reducedPartials_reducedPartials_sum_153 & partials_16_4; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_154 = reducedPartials_reducedPartials_carry_189 ^
    reducedPartials_reducedPartials_carry_188 ^ reducedPartials_reducedPartials_carry_187; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_190 = reducedPartials_reducedPartials_carry_189 &
    reducedPartials_reducedPartials_carry_188 | reducedPartials_reducedPartials_carry_188 &
    reducedPartials_reducedPartials_carry_187 | reducedPartials_reducedPartials_carry_189 &
    reducedPartials_reducedPartials_carry_187; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_155 = reducedPartials_reducedPartials_sum_154 ^
    reducedPartials_reducedPartials_carry_186 ^ partials_17_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_191 = reducedPartials_reducedPartials_sum_154 &
    reducedPartials_reducedPartials_carry_186 | reducedPartials_reducedPartials_carry_186 & partials_17_0 |
    reducedPartials_reducedPartials_sum_154 & partials_17_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_156 = reducedPartials_reducedPartials_sum_155 ^ partials_17_1 ^
    partials_17_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_192 = reducedPartials_reducedPartials_sum_155 & partials_17_1 |
    partials_17_1 & partials_17_2 | reducedPartials_reducedPartials_sum_155 & partials_17_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_157 = reducedPartials_reducedPartials_sum_156 ^ partials_17_3 ^
    partials_17_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_193 = reducedPartials_reducedPartials_sum_156 & partials_17_3 |
    partials_17_3 & partials_17_4 | reducedPartials_reducedPartials_sum_156 & partials_17_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_17_0 = reducedPartials_reducedPartials_sum_157 ^ partials_17_5; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_194 = reducedPartials_reducedPartials_sum_157 & partials_17_5; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_158 = reducedPartials_reducedPartials_carry_194 ^
    reducedPartials_reducedPartials_carry_193 ^ reducedPartials_reducedPartials_carry_192; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_195 = reducedPartials_reducedPartials_carry_194 &
    reducedPartials_reducedPartials_carry_193 | reducedPartials_reducedPartials_carry_193 &
    reducedPartials_reducedPartials_carry_192 | reducedPartials_reducedPartials_carry_194 &
    reducedPartials_reducedPartials_carry_192; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_159 = reducedPartials_reducedPartials_sum_158 ^
    reducedPartials_reducedPartials_carry_191 ^ reducedPartials_reducedPartials_carry_190; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_196 = reducedPartials_reducedPartials_sum_158 &
    reducedPartials_reducedPartials_carry_191 | reducedPartials_reducedPartials_carry_191 &
    reducedPartials_reducedPartials_carry_190 | reducedPartials_reducedPartials_sum_158 &
    reducedPartials_reducedPartials_carry_190; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_160 = reducedPartials_reducedPartials_sum_159 ^ partials_18_0 ^
    partials_18_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_197 = reducedPartials_reducedPartials_sum_159 & partials_18_0 |
    partials_18_0 & partials_18_1 | reducedPartials_reducedPartials_sum_159 & partials_18_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_161 = reducedPartials_reducedPartials_sum_160 ^ partials_18_2 ^
    partials_18_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_198 = reducedPartials_reducedPartials_sum_160 & partials_18_2 |
    partials_18_2 & partials_18_3 | reducedPartials_reducedPartials_sum_160 & partials_18_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_162 = reducedPartials_reducedPartials_sum_161 ^ partials_18_4 ^
    partials_18_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_199 = reducedPartials_reducedPartials_sum_161 & partials_18_4 |
    partials_18_4 & partials_18_5 | reducedPartials_reducedPartials_sum_161 & partials_18_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_18_0 = reducedPartials_reducedPartials_sum_162 ^ partials_18_6; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_200 = reducedPartials_reducedPartials_sum_162 & partials_18_6; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_163 = reducedPartials_reducedPartials_carry_200 ^
    reducedPartials_reducedPartials_carry_199 ^ reducedPartials_reducedPartials_carry_198; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_201 = reducedPartials_reducedPartials_carry_200 &
    reducedPartials_reducedPartials_carry_199 | reducedPartials_reducedPartials_carry_199 &
    reducedPartials_reducedPartials_carry_198 | reducedPartials_reducedPartials_carry_200 &
    reducedPartials_reducedPartials_carry_198; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_164 = reducedPartials_reducedPartials_sum_163 ^
    reducedPartials_reducedPartials_carry_197 ^ reducedPartials_reducedPartials_carry_196; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_202 = reducedPartials_reducedPartials_sum_163 &
    reducedPartials_reducedPartials_carry_197 | reducedPartials_reducedPartials_carry_197 &
    reducedPartials_reducedPartials_carry_196 | reducedPartials_reducedPartials_sum_163 &
    reducedPartials_reducedPartials_carry_196; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_165 = reducedPartials_reducedPartials_sum_164 ^
    reducedPartials_reducedPartials_carry_195 ^ reducedPartials_reducedPartials_19_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_203 = reducedPartials_reducedPartials_sum_164 &
    reducedPartials_reducedPartials_carry_195 | reducedPartials_reducedPartials_carry_195 &
    reducedPartials_reducedPartials_19_0 | reducedPartials_reducedPartials_sum_164 &
    reducedPartials_reducedPartials_19_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_166 = reducedPartials_reducedPartials_sum_165 ^ partials_19_2 ^
    partials_19_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_204 = reducedPartials_reducedPartials_sum_165 & partials_19_2 |
    partials_19_2 & partials_19_3 | reducedPartials_reducedPartials_sum_165 & partials_19_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_167 = reducedPartials_reducedPartials_sum_166 ^ partials_19_4 ^
    partials_19_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_205 = reducedPartials_reducedPartials_sum_166 & partials_19_4 |
    partials_19_4 & partials_19_5 | reducedPartials_reducedPartials_sum_166 & partials_19_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_19_0_1 = reducedPartials_reducedPartials_sum_167 ^ partials_19_6 ^ partials_19_7
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_206 = reducedPartials_reducedPartials_sum_167 & partials_19_6 |
    partials_19_6 & partials_19_7 | reducedPartials_reducedPartials_sum_167 & partials_19_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_168 = reducedPartials_reducedPartials_carry_206 ^
    reducedPartials_reducedPartials_carry_205 ^ reducedPartials_reducedPartials_carry_204; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_207 = reducedPartials_reducedPartials_carry_206 &
    reducedPartials_reducedPartials_carry_205 | reducedPartials_reducedPartials_carry_205 &
    reducedPartials_reducedPartials_carry_204 | reducedPartials_reducedPartials_carry_206 &
    reducedPartials_reducedPartials_carry_204; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_169 = reducedPartials_reducedPartials_sum_168 ^
    reducedPartials_reducedPartials_carry_203 ^ reducedPartials_reducedPartials_carry_202; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_208 = reducedPartials_reducedPartials_sum_168 &
    reducedPartials_reducedPartials_carry_203 | reducedPartials_reducedPartials_carry_203 &
    reducedPartials_reducedPartials_carry_202 | reducedPartials_reducedPartials_sum_168 &
    reducedPartials_reducedPartials_carry_202; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_170 = reducedPartials_reducedPartials_sum_169 ^
    reducedPartials_reducedPartials_carry_201 ^ reducedPartials_reducedPartials_20_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_209 = reducedPartials_reducedPartials_sum_169 &
    reducedPartials_reducedPartials_carry_201 | reducedPartials_reducedPartials_carry_201 &
    reducedPartials_reducedPartials_20_0 | reducedPartials_reducedPartials_sum_169 &
    reducedPartials_reducedPartials_20_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_171 = reducedPartials_reducedPartials_sum_170 ^ partials_20_3 ^
    partials_20_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_210 = reducedPartials_reducedPartials_sum_170 & partials_20_3 |
    partials_20_3 & partials_20_4 | reducedPartials_reducedPartials_sum_170 & partials_20_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_172 = reducedPartials_reducedPartials_sum_171 ^ partials_20_5 ^
    partials_20_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_211 = reducedPartials_reducedPartials_sum_171 & partials_20_5 |
    partials_20_5 & partials_20_6 | reducedPartials_reducedPartials_sum_171 & partials_20_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_20_0_1 = reducedPartials_reducedPartials_sum_172 ^ partials_20_7 ^ partials_20_8
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_212 = reducedPartials_reducedPartials_sum_172 & partials_20_7 |
    partials_20_7 & partials_20_8 | reducedPartials_reducedPartials_sum_172 & partials_20_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_173 = reducedPartials_reducedPartials_carry_212 ^
    reducedPartials_reducedPartials_carry_211 ^ reducedPartials_reducedPartials_carry_210; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_213 = reducedPartials_reducedPartials_carry_212 &
    reducedPartials_reducedPartials_carry_211 | reducedPartials_reducedPartials_carry_211 &
    reducedPartials_reducedPartials_carry_210 | reducedPartials_reducedPartials_carry_212 &
    reducedPartials_reducedPartials_carry_210; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_174 = reducedPartials_reducedPartials_sum_173 ^
    reducedPartials_reducedPartials_carry_209 ^ reducedPartials_reducedPartials_carry_208; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_214 = reducedPartials_reducedPartials_sum_173 &
    reducedPartials_reducedPartials_carry_209 | reducedPartials_reducedPartials_carry_209 &
    reducedPartials_reducedPartials_carry_208 | reducedPartials_reducedPartials_sum_173 &
    reducedPartials_reducedPartials_carry_208; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_175 = reducedPartials_reducedPartials_sum_174 ^
    reducedPartials_reducedPartials_carry_207 ^ reducedPartials_reducedPartials_21_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_215 = reducedPartials_reducedPartials_sum_174 &
    reducedPartials_reducedPartials_carry_207 | reducedPartials_reducedPartials_carry_207 &
    reducedPartials_reducedPartials_21_0 | reducedPartials_reducedPartials_sum_174 &
    reducedPartials_reducedPartials_21_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_176 = reducedPartials_reducedPartials_sum_175 ^ partials_21_4 ^
    partials_21_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_216 = reducedPartials_reducedPartials_sum_175 & partials_21_4 |
    partials_21_4 & partials_21_5 | reducedPartials_reducedPartials_sum_175 & partials_21_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_177 = reducedPartials_reducedPartials_sum_176 ^ partials_21_6 ^
    partials_21_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_217 = reducedPartials_reducedPartials_sum_176 & partials_21_6 |
    partials_21_6 & partials_21_7 | reducedPartials_reducedPartials_sum_176 & partials_21_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_21_0_1 = reducedPartials_reducedPartials_sum_177 ^ partials_21_8 ^ partials_21_9
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_218 = reducedPartials_reducedPartials_sum_177 & partials_21_8 |
    partials_21_8 & partials_21_9 | reducedPartials_reducedPartials_sum_177 & partials_21_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_178 = reducedPartials_reducedPartials_carry_218 ^
    reducedPartials_reducedPartials_carry_217 ^ reducedPartials_reducedPartials_carry_216; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_219 = reducedPartials_reducedPartials_carry_218 &
    reducedPartials_reducedPartials_carry_217 | reducedPartials_reducedPartials_carry_217 &
    reducedPartials_reducedPartials_carry_216 | reducedPartials_reducedPartials_carry_218 &
    reducedPartials_reducedPartials_carry_216; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_179 = reducedPartials_reducedPartials_sum_178 ^
    reducedPartials_reducedPartials_carry_215 ^ reducedPartials_reducedPartials_carry_214; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_220 = reducedPartials_reducedPartials_sum_178 &
    reducedPartials_reducedPartials_carry_215 | reducedPartials_reducedPartials_carry_215 &
    reducedPartials_reducedPartials_carry_214 | reducedPartials_reducedPartials_sum_178 &
    reducedPartials_reducedPartials_carry_214; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_180 = reducedPartials_reducedPartials_sum_179 ^
    reducedPartials_reducedPartials_carry_213 ^ reducedPartials_reducedPartials_22_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_221 = reducedPartials_reducedPartials_sum_179 &
    reducedPartials_reducedPartials_carry_213 | reducedPartials_reducedPartials_carry_213 &
    reducedPartials_reducedPartials_22_0 | reducedPartials_reducedPartials_sum_179 &
    reducedPartials_reducedPartials_22_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_181 = reducedPartials_reducedPartials_sum_180 ^ partials_22_5 ^
    partials_22_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_222 = reducedPartials_reducedPartials_sum_180 & partials_22_5 |
    partials_22_5 & partials_22_6 | reducedPartials_reducedPartials_sum_180 & partials_22_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_182 = reducedPartials_reducedPartials_sum_181 ^ partials_22_7 ^
    partials_22_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_223 = reducedPartials_reducedPartials_sum_181 & partials_22_7 |
    partials_22_7 & partials_22_8 | reducedPartials_reducedPartials_sum_181 & partials_22_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_22_0_1 = reducedPartials_reducedPartials_sum_182 ^ partials_22_9 ^
    partials_22_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_224 = reducedPartials_reducedPartials_sum_182 & partials_22_9 |
    partials_22_9 & partials_22_10 | reducedPartials_reducedPartials_sum_182 & partials_22_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_183 = reducedPartials_reducedPartials_carry_224 ^
    reducedPartials_reducedPartials_carry_223 ^ reducedPartials_reducedPartials_carry_222; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_225 = reducedPartials_reducedPartials_carry_224 &
    reducedPartials_reducedPartials_carry_223 | reducedPartials_reducedPartials_carry_223 &
    reducedPartials_reducedPartials_carry_222 | reducedPartials_reducedPartials_carry_224 &
    reducedPartials_reducedPartials_carry_222; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_184 = reducedPartials_reducedPartials_sum_183 ^
    reducedPartials_reducedPartials_carry_221 ^ reducedPartials_reducedPartials_carry_220; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_226 = reducedPartials_reducedPartials_sum_183 &
    reducedPartials_reducedPartials_carry_221 | reducedPartials_reducedPartials_carry_221 &
    reducedPartials_reducedPartials_carry_220 | reducedPartials_reducedPartials_sum_183 &
    reducedPartials_reducedPartials_carry_220; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_185 = reducedPartials_reducedPartials_sum_184 ^
    reducedPartials_reducedPartials_carry_219 ^ reducedPartials_reducedPartials_23_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_227 = reducedPartials_reducedPartials_sum_184 &
    reducedPartials_reducedPartials_carry_219 | reducedPartials_reducedPartials_carry_219 &
    reducedPartials_reducedPartials_23_0 | reducedPartials_reducedPartials_sum_184 &
    reducedPartials_reducedPartials_23_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_186 = reducedPartials_reducedPartials_sum_185 ^ partials_23_6 ^
    partials_23_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_228 = reducedPartials_reducedPartials_sum_185 & partials_23_6 |
    partials_23_6 & partials_23_7 | reducedPartials_reducedPartials_sum_185 & partials_23_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_187 = reducedPartials_reducedPartials_sum_186 ^ partials_23_8 ^
    partials_23_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_229 = reducedPartials_reducedPartials_sum_186 & partials_23_8 |
    partials_23_8 & partials_23_9 | reducedPartials_reducedPartials_sum_186 & partials_23_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_23_0_1 = reducedPartials_reducedPartials_sum_187 ^ partials_23_10 ^
    partials_23_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_230 = reducedPartials_reducedPartials_sum_187 & partials_23_10 |
    partials_23_10 & partials_23_11 | reducedPartials_reducedPartials_sum_187 & partials_23_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_188 = reducedPartials_reducedPartials_carry_230 ^
    reducedPartials_reducedPartials_carry_229 ^ reducedPartials_reducedPartials_carry_228; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_231 = reducedPartials_reducedPartials_carry_230 &
    reducedPartials_reducedPartials_carry_229 | reducedPartials_reducedPartials_carry_229 &
    reducedPartials_reducedPartials_carry_228 | reducedPartials_reducedPartials_carry_230 &
    reducedPartials_reducedPartials_carry_228; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_189 = reducedPartials_reducedPartials_sum_188 ^
    reducedPartials_reducedPartials_carry_227 ^ reducedPartials_reducedPartials_carry_226; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_232 = reducedPartials_reducedPartials_sum_188 &
    reducedPartials_reducedPartials_carry_227 | reducedPartials_reducedPartials_carry_227 &
    reducedPartials_reducedPartials_carry_226 | reducedPartials_reducedPartials_sum_188 &
    reducedPartials_reducedPartials_carry_226; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_190 = reducedPartials_reducedPartials_sum_189 ^
    reducedPartials_reducedPartials_carry_225 ^ reducedPartials_reducedPartials_24_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_233 = reducedPartials_reducedPartials_sum_189 &
    reducedPartials_reducedPartials_carry_225 | reducedPartials_reducedPartials_carry_225 &
    reducedPartials_reducedPartials_24_0 | reducedPartials_reducedPartials_sum_189 &
    reducedPartials_reducedPartials_24_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_191 = reducedPartials_reducedPartials_sum_190 ^ partials_24_7 ^
    partials_24_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_234 = reducedPartials_reducedPartials_sum_190 & partials_24_7 |
    partials_24_7 & partials_24_8 | reducedPartials_reducedPartials_sum_190 & partials_24_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_192 = reducedPartials_reducedPartials_sum_191 ^ partials_24_9 ^
    partials_24_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_235 = reducedPartials_reducedPartials_sum_191 & partials_24_9 |
    partials_24_9 & partials_24_10 | reducedPartials_reducedPartials_sum_191 & partials_24_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_24_0_1 = reducedPartials_reducedPartials_sum_192 ^ partials_24_11 ^
    partials_24_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_236 = reducedPartials_reducedPartials_sum_192 & partials_24_11 |
    partials_24_11 & partials_24_12 | reducedPartials_reducedPartials_sum_192 & partials_24_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_193 = reducedPartials_reducedPartials_carry_236 ^
    reducedPartials_reducedPartials_carry_235 ^ reducedPartials_reducedPartials_carry_234; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_237 = reducedPartials_reducedPartials_carry_236 &
    reducedPartials_reducedPartials_carry_235 | reducedPartials_reducedPartials_carry_235 &
    reducedPartials_reducedPartials_carry_234 | reducedPartials_reducedPartials_carry_236 &
    reducedPartials_reducedPartials_carry_234; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_194 = reducedPartials_reducedPartials_sum_193 ^
    reducedPartials_reducedPartials_carry_233 ^ reducedPartials_reducedPartials_carry_232; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_238 = reducedPartials_reducedPartials_sum_193 &
    reducedPartials_reducedPartials_carry_233 | reducedPartials_reducedPartials_carry_233 &
    reducedPartials_reducedPartials_carry_232 | reducedPartials_reducedPartials_sum_193 &
    reducedPartials_reducedPartials_carry_232; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_195 = reducedPartials_reducedPartials_sum_194 ^
    reducedPartials_reducedPartials_carry_231 ^ reducedPartials_reducedPartials_25_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_239 = reducedPartials_reducedPartials_sum_194 &
    reducedPartials_reducedPartials_carry_231 | reducedPartials_reducedPartials_carry_231 &
    reducedPartials_reducedPartials_25_0 | reducedPartials_reducedPartials_sum_194 &
    reducedPartials_reducedPartials_25_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_196 = reducedPartials_reducedPartials_sum_195 ^ partials_25_8 ^
    partials_25_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_240 = reducedPartials_reducedPartials_sum_195 & partials_25_8 |
    partials_25_8 & partials_25_9 | reducedPartials_reducedPartials_sum_195 & partials_25_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_197 = reducedPartials_reducedPartials_sum_196 ^ partials_25_10 ^
    partials_25_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_241 = reducedPartials_reducedPartials_sum_196 & partials_25_10 |
    partials_25_10 & partials_25_11 | reducedPartials_reducedPartials_sum_196 & partials_25_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_25_0_1 = reducedPartials_reducedPartials_sum_197 ^ partials_25_12 ^
    partials_25_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_242 = reducedPartials_reducedPartials_sum_197 & partials_25_12 |
    partials_25_12 & partials_25_13 | reducedPartials_reducedPartials_sum_197 & partials_25_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_198 = reducedPartials_reducedPartials_carry_242 ^
    reducedPartials_reducedPartials_carry_241 ^ reducedPartials_reducedPartials_carry_240; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_243 = reducedPartials_reducedPartials_carry_242 &
    reducedPartials_reducedPartials_carry_241 | reducedPartials_reducedPartials_carry_241 &
    reducedPartials_reducedPartials_carry_240 | reducedPartials_reducedPartials_carry_242 &
    reducedPartials_reducedPartials_carry_240; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_199 = reducedPartials_reducedPartials_sum_198 ^
    reducedPartials_reducedPartials_carry_239 ^ reducedPartials_reducedPartials_carry_238; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_244 = reducedPartials_reducedPartials_sum_198 &
    reducedPartials_reducedPartials_carry_239 | reducedPartials_reducedPartials_carry_239 &
    reducedPartials_reducedPartials_carry_238 | reducedPartials_reducedPartials_sum_198 &
    reducedPartials_reducedPartials_carry_238; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_200 = reducedPartials_reducedPartials_sum_199 ^
    reducedPartials_reducedPartials_carry_237 ^ reducedPartials_reducedPartials_26_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_245 = reducedPartials_reducedPartials_sum_199 &
    reducedPartials_reducedPartials_carry_237 | reducedPartials_reducedPartials_carry_237 &
    reducedPartials_reducedPartials_26_0 | reducedPartials_reducedPartials_sum_199 &
    reducedPartials_reducedPartials_26_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_201 = reducedPartials_reducedPartials_sum_200 ^ partials_26_9 ^
    partials_26_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_246 = reducedPartials_reducedPartials_sum_200 & partials_26_9 |
    partials_26_9 & partials_26_10 | reducedPartials_reducedPartials_sum_200 & partials_26_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_202 = reducedPartials_reducedPartials_sum_201 ^ partials_26_11 ^
    partials_26_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_247 = reducedPartials_reducedPartials_sum_201 & partials_26_11 |
    partials_26_11 & partials_26_12 | reducedPartials_reducedPartials_sum_201 & partials_26_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_26_0_1 = reducedPartials_reducedPartials_sum_202 ^ partials_26_13 ^
    partials_26_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_248 = reducedPartials_reducedPartials_sum_202 & partials_26_13 |
    partials_26_13 & partials_26_14 | reducedPartials_reducedPartials_sum_202 & partials_26_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_203 = reducedPartials_reducedPartials_carry_248 ^
    reducedPartials_reducedPartials_carry_247 ^ reducedPartials_reducedPartials_carry_246; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_249 = reducedPartials_reducedPartials_carry_248 &
    reducedPartials_reducedPartials_carry_247 | reducedPartials_reducedPartials_carry_247 &
    reducedPartials_reducedPartials_carry_246 | reducedPartials_reducedPartials_carry_248 &
    reducedPartials_reducedPartials_carry_246; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_204 = reducedPartials_reducedPartials_sum_203 ^
    reducedPartials_reducedPartials_carry_245 ^ reducedPartials_reducedPartials_carry_244; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_250 = reducedPartials_reducedPartials_sum_203 &
    reducedPartials_reducedPartials_carry_245 | reducedPartials_reducedPartials_carry_245 &
    reducedPartials_reducedPartials_carry_244 | reducedPartials_reducedPartials_sum_203 &
    reducedPartials_reducedPartials_carry_244; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_205 = reducedPartials_reducedPartials_sum_204 ^
    reducedPartials_reducedPartials_carry_243 ^ reducedPartials_reducedPartials_27_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_251 = reducedPartials_reducedPartials_sum_204 &
    reducedPartials_reducedPartials_carry_243 | reducedPartials_reducedPartials_carry_243 &
    reducedPartials_reducedPartials_27_0 | reducedPartials_reducedPartials_sum_204 &
    reducedPartials_reducedPartials_27_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_206 = reducedPartials_reducedPartials_sum_205 ^ partials_27_10 ^
    partials_27_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_252 = reducedPartials_reducedPartials_sum_205 & partials_27_10 |
    partials_27_10 & partials_27_11 | reducedPartials_reducedPartials_sum_205 & partials_27_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_207 = reducedPartials_reducedPartials_sum_206 ^ partials_27_12 ^
    partials_27_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_253 = reducedPartials_reducedPartials_sum_206 & partials_27_12 |
    partials_27_12 & partials_27_13 | reducedPartials_reducedPartials_sum_206 & partials_27_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_27_0_1 = reducedPartials_reducedPartials_sum_207 ^ partials_27_14 ^
    partials_27_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_254 = reducedPartials_reducedPartials_sum_207 & partials_27_14 |
    partials_27_14 & partials_27_15 | reducedPartials_reducedPartials_sum_207 & partials_27_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_208 = reducedPartials_reducedPartials_carry_254 ^
    reducedPartials_reducedPartials_carry_253 ^ reducedPartials_reducedPartials_carry_252; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_255 = reducedPartials_reducedPartials_carry_254 &
    reducedPartials_reducedPartials_carry_253 | reducedPartials_reducedPartials_carry_253 &
    reducedPartials_reducedPartials_carry_252 | reducedPartials_reducedPartials_carry_254 &
    reducedPartials_reducedPartials_carry_252; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_209 = reducedPartials_reducedPartials_sum_208 ^
    reducedPartials_reducedPartials_carry_251 ^ reducedPartials_reducedPartials_carry_250; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_256 = reducedPartials_reducedPartials_sum_208 &
    reducedPartials_reducedPartials_carry_251 | reducedPartials_reducedPartials_carry_251 &
    reducedPartials_reducedPartials_carry_250 | reducedPartials_reducedPartials_sum_208 &
    reducedPartials_reducedPartials_carry_250; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_210 = reducedPartials_reducedPartials_sum_209 ^
    reducedPartials_reducedPartials_carry_249 ^ reducedPartials_reducedPartials_28_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_257 = reducedPartials_reducedPartials_sum_209 &
    reducedPartials_reducedPartials_carry_249 | reducedPartials_reducedPartials_carry_249 &
    reducedPartials_reducedPartials_28_0_1 | reducedPartials_reducedPartials_sum_209 &
    reducedPartials_reducedPartials_28_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_211 = reducedPartials_reducedPartials_sum_210 ^ partials_28_11 ^
    partials_28_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_258 = reducedPartials_reducedPartials_sum_210 & partials_28_11 |
    partials_28_11 & partials_28_12 | reducedPartials_reducedPartials_sum_210 & partials_28_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_212 = reducedPartials_reducedPartials_sum_211 ^ partials_28_13 ^
    partials_28_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_259 = reducedPartials_reducedPartials_sum_211 & partials_28_13 |
    partials_28_13 & partials_28_14 | reducedPartials_reducedPartials_sum_211 & partials_28_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_28_0_2 = reducedPartials_reducedPartials_sum_212 ^ partials_28_15 ^
    partials_28_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_260 = reducedPartials_reducedPartials_sum_212 & partials_28_15 |
    partials_28_15 & partials_28_16 | reducedPartials_reducedPartials_sum_212 & partials_28_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_213 = reducedPartials_reducedPartials_carry_260 ^
    reducedPartials_reducedPartials_carry_259 ^ reducedPartials_reducedPartials_carry_258; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_261 = reducedPartials_reducedPartials_carry_260 &
    reducedPartials_reducedPartials_carry_259 | reducedPartials_reducedPartials_carry_259 &
    reducedPartials_reducedPartials_carry_258 | reducedPartials_reducedPartials_carry_260 &
    reducedPartials_reducedPartials_carry_258; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_214 = reducedPartials_reducedPartials_sum_213 ^
    reducedPartials_reducedPartials_carry_257 ^ reducedPartials_reducedPartials_carry_256; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_262 = reducedPartials_reducedPartials_sum_213 &
    reducedPartials_reducedPartials_carry_257 | reducedPartials_reducedPartials_carry_257 &
    reducedPartials_reducedPartials_carry_256 | reducedPartials_reducedPartials_sum_213 &
    reducedPartials_reducedPartials_carry_256; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_215 = reducedPartials_reducedPartials_sum_214 ^
    reducedPartials_reducedPartials_carry_255 ^ reducedPartials_reducedPartials_29_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_263 = reducedPartials_reducedPartials_sum_214 &
    reducedPartials_reducedPartials_carry_255 | reducedPartials_reducedPartials_carry_255 &
    reducedPartials_reducedPartials_29_0_1 | reducedPartials_reducedPartials_sum_214 &
    reducedPartials_reducedPartials_29_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_216 = reducedPartials_reducedPartials_sum_215 ^ partials_29_12 ^
    partials_29_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_264 = reducedPartials_reducedPartials_sum_215 & partials_29_12 |
    partials_29_12 & partials_29_13 | reducedPartials_reducedPartials_sum_215 & partials_29_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_217 = reducedPartials_reducedPartials_sum_216 ^ partials_29_14 ^
    partials_29_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_265 = reducedPartials_reducedPartials_sum_216 & partials_29_14 |
    partials_29_14 & partials_29_15 | reducedPartials_reducedPartials_sum_216 & partials_29_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_29_0_2 = reducedPartials_reducedPartials_sum_217 ^ partials_29_16 ^
    partials_29_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_266 = reducedPartials_reducedPartials_sum_217 & partials_29_16 |
    partials_29_16 & partials_29_17 | reducedPartials_reducedPartials_sum_217 & partials_29_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_218 = reducedPartials_reducedPartials_carry_266 ^
    reducedPartials_reducedPartials_carry_265 ^ reducedPartials_reducedPartials_carry_264; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_267 = reducedPartials_reducedPartials_carry_266 &
    reducedPartials_reducedPartials_carry_265 | reducedPartials_reducedPartials_carry_265 &
    reducedPartials_reducedPartials_carry_264 | reducedPartials_reducedPartials_carry_266 &
    reducedPartials_reducedPartials_carry_264; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_219 = reducedPartials_reducedPartials_sum_218 ^
    reducedPartials_reducedPartials_carry_263 ^ reducedPartials_reducedPartials_carry_262; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_268 = reducedPartials_reducedPartials_sum_218 &
    reducedPartials_reducedPartials_carry_263 | reducedPartials_reducedPartials_carry_263 &
    reducedPartials_reducedPartials_carry_262 | reducedPartials_reducedPartials_sum_218 &
    reducedPartials_reducedPartials_carry_262; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_220 = reducedPartials_reducedPartials_sum_219 ^
    reducedPartials_reducedPartials_carry_261 ^ reducedPartials_reducedPartials_30_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_269 = reducedPartials_reducedPartials_sum_219 &
    reducedPartials_reducedPartials_carry_261 | reducedPartials_reducedPartials_carry_261 &
    reducedPartials_reducedPartials_30_0_1 | reducedPartials_reducedPartials_sum_219 &
    reducedPartials_reducedPartials_30_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_221 = reducedPartials_reducedPartials_sum_220 ^ partials_30_13 ^
    partials_30_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_270 = reducedPartials_reducedPartials_sum_220 & partials_30_13 |
    partials_30_13 & partials_30_14 | reducedPartials_reducedPartials_sum_220 & partials_30_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_222 = reducedPartials_reducedPartials_sum_221 ^ partials_30_15 ^
    partials_30_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_271 = reducedPartials_reducedPartials_sum_221 & partials_30_15 |
    partials_30_15 & partials_30_16 | reducedPartials_reducedPartials_sum_221 & partials_30_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_30_0_2 = reducedPartials_reducedPartials_sum_222 ^ partials_30_17 ^
    partials_30_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_272 = reducedPartials_reducedPartials_sum_222 & partials_30_17 |
    partials_30_17 & partials_30_18 | reducedPartials_reducedPartials_sum_222 & partials_30_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_223 = reducedPartials_reducedPartials_carry_272 ^
    reducedPartials_reducedPartials_carry_271 ^ reducedPartials_reducedPartials_carry_270; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_273 = reducedPartials_reducedPartials_carry_272 &
    reducedPartials_reducedPartials_carry_271 | reducedPartials_reducedPartials_carry_271 &
    reducedPartials_reducedPartials_carry_270 | reducedPartials_reducedPartials_carry_272 &
    reducedPartials_reducedPartials_carry_270; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_224 = reducedPartials_reducedPartials_sum_223 ^
    reducedPartials_reducedPartials_carry_269 ^ reducedPartials_reducedPartials_carry_268; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_274 = reducedPartials_reducedPartials_sum_223 &
    reducedPartials_reducedPartials_carry_269 | reducedPartials_reducedPartials_carry_269 &
    reducedPartials_reducedPartials_carry_268 | reducedPartials_reducedPartials_sum_223 &
    reducedPartials_reducedPartials_carry_268; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_225 = reducedPartials_reducedPartials_sum_224 ^
    reducedPartials_reducedPartials_carry_267 ^ reducedPartials_reducedPartials_31_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_275 = reducedPartials_reducedPartials_sum_224 &
    reducedPartials_reducedPartials_carry_267 | reducedPartials_reducedPartials_carry_267 &
    reducedPartials_reducedPartials_31_0_1 | reducedPartials_reducedPartials_sum_224 &
    reducedPartials_reducedPartials_31_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_226 = reducedPartials_reducedPartials_sum_225 ^ partials_31_14 ^
    partials_31_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_276 = reducedPartials_reducedPartials_sum_225 & partials_31_14 |
    partials_31_14 & partials_31_15 | reducedPartials_reducedPartials_sum_225 & partials_31_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_227 = reducedPartials_reducedPartials_sum_226 ^ partials_31_16 ^
    partials_31_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_277 = reducedPartials_reducedPartials_sum_226 & partials_31_16 |
    partials_31_16 & partials_31_17 | reducedPartials_reducedPartials_sum_226 & partials_31_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_31_0_2 = reducedPartials_reducedPartials_sum_227 ^ partials_31_18 ^
    partials_31_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_278 = reducedPartials_reducedPartials_sum_227 & partials_31_18 |
    partials_31_18 & partials_31_19 | reducedPartials_reducedPartials_sum_227 & partials_31_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_228 = reducedPartials_reducedPartials_carry_278 ^
    reducedPartials_reducedPartials_carry_277 ^ reducedPartials_reducedPartials_carry_276; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_279 = reducedPartials_reducedPartials_carry_278 &
    reducedPartials_reducedPartials_carry_277 | reducedPartials_reducedPartials_carry_277 &
    reducedPartials_reducedPartials_carry_276 | reducedPartials_reducedPartials_carry_278 &
    reducedPartials_reducedPartials_carry_276; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_229 = reducedPartials_reducedPartials_sum_228 ^
    reducedPartials_reducedPartials_carry_275 ^ reducedPartials_reducedPartials_carry_274; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_280 = reducedPartials_reducedPartials_sum_228 &
    reducedPartials_reducedPartials_carry_275 | reducedPartials_reducedPartials_carry_275 &
    reducedPartials_reducedPartials_carry_274 | reducedPartials_reducedPartials_sum_228 &
    reducedPartials_reducedPartials_carry_274; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_230 = reducedPartials_reducedPartials_sum_229 ^
    reducedPartials_reducedPartials_carry_273 ^ reducedPartials_reducedPartials_32_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_281 = reducedPartials_reducedPartials_sum_229 &
    reducedPartials_reducedPartials_carry_273 | reducedPartials_reducedPartials_carry_273 &
    reducedPartials_reducedPartials_32_0_1 | reducedPartials_reducedPartials_sum_229 &
    reducedPartials_reducedPartials_32_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_231 = reducedPartials_reducedPartials_sum_230 ^ partials_32_13 ^
    partials_32_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_282 = reducedPartials_reducedPartials_sum_230 & partials_32_13 |
    partials_32_13 & partials_32_14 | reducedPartials_reducedPartials_sum_230 & partials_32_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_232 = reducedPartials_reducedPartials_sum_231 ^ partials_32_15 ^
    partials_32_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_283 = reducedPartials_reducedPartials_sum_231 & partials_32_15 |
    partials_32_15 & partials_32_16 | reducedPartials_reducedPartials_sum_231 & partials_32_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_32_0_2 = reducedPartials_reducedPartials_sum_232 ^ partials_32_17 ^
    partials_32_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_284 = reducedPartials_reducedPartials_sum_232 & partials_32_17 |
    partials_32_17 & partials_32_18 | reducedPartials_reducedPartials_sum_232 & partials_32_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_233 = reducedPartials_reducedPartials_carry_284 ^
    reducedPartials_reducedPartials_carry_283 ^ reducedPartials_reducedPartials_carry_282; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_285 = reducedPartials_reducedPartials_carry_284 &
    reducedPartials_reducedPartials_carry_283 | reducedPartials_reducedPartials_carry_283 &
    reducedPartials_reducedPartials_carry_282 | reducedPartials_reducedPartials_carry_284 &
    reducedPartials_reducedPartials_carry_282; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_234 = reducedPartials_reducedPartials_sum_233 ^
    reducedPartials_reducedPartials_carry_281 ^ reducedPartials_reducedPartials_carry_280; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_286 = reducedPartials_reducedPartials_sum_233 &
    reducedPartials_reducedPartials_carry_281 | reducedPartials_reducedPartials_carry_281 &
    reducedPartials_reducedPartials_carry_280 | reducedPartials_reducedPartials_sum_233 &
    reducedPartials_reducedPartials_carry_280; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_235 = reducedPartials_reducedPartials_sum_234 ^
    reducedPartials_reducedPartials_carry_279 ^ reducedPartials_reducedPartials_33_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_287 = reducedPartials_reducedPartials_sum_234 &
    reducedPartials_reducedPartials_carry_279 | reducedPartials_reducedPartials_carry_279 &
    reducedPartials_reducedPartials_33_0_1 | reducedPartials_reducedPartials_sum_234 &
    reducedPartials_reducedPartials_33_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_236 = reducedPartials_reducedPartials_sum_235 ^ partials_33_12 ^
    partials_33_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_288 = reducedPartials_reducedPartials_sum_235 & partials_33_12 |
    partials_33_12 & partials_33_13 | reducedPartials_reducedPartials_sum_235 & partials_33_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_237 = reducedPartials_reducedPartials_sum_236 ^ partials_33_14 ^
    partials_33_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_289 = reducedPartials_reducedPartials_sum_236 & partials_33_14 |
    partials_33_14 & partials_33_15 | reducedPartials_reducedPartials_sum_236 & partials_33_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_33_0_2 = reducedPartials_reducedPartials_sum_237 ^ partials_33_16 ^
    partials_33_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_290 = reducedPartials_reducedPartials_sum_237 & partials_33_16 |
    partials_33_16 & partials_33_17 | reducedPartials_reducedPartials_sum_237 & partials_33_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_238 = reducedPartials_reducedPartials_carry_290 ^
    reducedPartials_reducedPartials_carry_289 ^ reducedPartials_reducedPartials_carry_288; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_291 = reducedPartials_reducedPartials_carry_290 &
    reducedPartials_reducedPartials_carry_289 | reducedPartials_reducedPartials_carry_289 &
    reducedPartials_reducedPartials_carry_288 | reducedPartials_reducedPartials_carry_290 &
    reducedPartials_reducedPartials_carry_288; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_239 = reducedPartials_reducedPartials_sum_238 ^
    reducedPartials_reducedPartials_carry_287 ^ reducedPartials_reducedPartials_carry_286; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_292 = reducedPartials_reducedPartials_sum_238 &
    reducedPartials_reducedPartials_carry_287 | reducedPartials_reducedPartials_carry_287 &
    reducedPartials_reducedPartials_carry_286 | reducedPartials_reducedPartials_sum_238 &
    reducedPartials_reducedPartials_carry_286; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_240 = reducedPartials_reducedPartials_sum_239 ^
    reducedPartials_reducedPartials_carry_285 ^ reducedPartials_reducedPartials_34_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_293 = reducedPartials_reducedPartials_sum_239 &
    reducedPartials_reducedPartials_carry_285 | reducedPartials_reducedPartials_carry_285 &
    reducedPartials_reducedPartials_34_0_1 | reducedPartials_reducedPartials_sum_239 &
    reducedPartials_reducedPartials_34_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_241 = reducedPartials_reducedPartials_sum_240 ^ partials_34_11 ^
    partials_34_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_294 = reducedPartials_reducedPartials_sum_240 & partials_34_11 |
    partials_34_11 & partials_34_12 | reducedPartials_reducedPartials_sum_240 & partials_34_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_242 = reducedPartials_reducedPartials_sum_241 ^ partials_34_13 ^
    partials_34_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_295 = reducedPartials_reducedPartials_sum_241 & partials_34_13 |
    partials_34_13 & partials_34_14 | reducedPartials_reducedPartials_sum_241 & partials_34_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_34_0_2 = reducedPartials_reducedPartials_sum_242 ^ partials_34_15 ^
    partials_34_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_296 = reducedPartials_reducedPartials_sum_242 & partials_34_15 |
    partials_34_15 & partials_34_16 | reducedPartials_reducedPartials_sum_242 & partials_34_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_243 = reducedPartials_reducedPartials_carry_296 ^
    reducedPartials_reducedPartials_carry_295 ^ reducedPartials_reducedPartials_carry_294; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_297 = reducedPartials_reducedPartials_carry_296 &
    reducedPartials_reducedPartials_carry_295 | reducedPartials_reducedPartials_carry_295 &
    reducedPartials_reducedPartials_carry_294 | reducedPartials_reducedPartials_carry_296 &
    reducedPartials_reducedPartials_carry_294; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_244 = reducedPartials_reducedPartials_sum_243 ^
    reducedPartials_reducedPartials_carry_293 ^ reducedPartials_reducedPartials_carry_292; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_298 = reducedPartials_reducedPartials_sum_243 &
    reducedPartials_reducedPartials_carry_293 | reducedPartials_reducedPartials_carry_293 &
    reducedPartials_reducedPartials_carry_292 | reducedPartials_reducedPartials_sum_243 &
    reducedPartials_reducedPartials_carry_292; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_245 = reducedPartials_reducedPartials_sum_244 ^
    reducedPartials_reducedPartials_carry_291 ^ reducedPartials_reducedPartials_35_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_299 = reducedPartials_reducedPartials_sum_244 &
    reducedPartials_reducedPartials_carry_291 | reducedPartials_reducedPartials_carry_291 &
    reducedPartials_reducedPartials_35_0_1 | reducedPartials_reducedPartials_sum_244 &
    reducedPartials_reducedPartials_35_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_246 = reducedPartials_reducedPartials_sum_245 ^ partials_35_10 ^
    partials_35_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_300 = reducedPartials_reducedPartials_sum_245 & partials_35_10 |
    partials_35_10 & partials_35_11 | reducedPartials_reducedPartials_sum_245 & partials_35_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_247 = reducedPartials_reducedPartials_sum_246 ^ partials_35_12 ^
    partials_35_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_301 = reducedPartials_reducedPartials_sum_246 & partials_35_12 |
    partials_35_12 & partials_35_13 | reducedPartials_reducedPartials_sum_246 & partials_35_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_35_0_2 = reducedPartials_reducedPartials_sum_247 ^ partials_35_14 ^
    partials_35_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_302 = reducedPartials_reducedPartials_sum_247 & partials_35_14 |
    partials_35_14 & partials_35_15 | reducedPartials_reducedPartials_sum_247 & partials_35_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_248 = reducedPartials_reducedPartials_carry_302 ^
    reducedPartials_reducedPartials_carry_301 ^ reducedPartials_reducedPartials_carry_300; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_303 = reducedPartials_reducedPartials_carry_302 &
    reducedPartials_reducedPartials_carry_301 | reducedPartials_reducedPartials_carry_301 &
    reducedPartials_reducedPartials_carry_300 | reducedPartials_reducedPartials_carry_302 &
    reducedPartials_reducedPartials_carry_300; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_249 = reducedPartials_reducedPartials_sum_248 ^
    reducedPartials_reducedPartials_carry_299 ^ reducedPartials_reducedPartials_carry_298; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_304 = reducedPartials_reducedPartials_sum_248 &
    reducedPartials_reducedPartials_carry_299 | reducedPartials_reducedPartials_carry_299 &
    reducedPartials_reducedPartials_carry_298 | reducedPartials_reducedPartials_sum_248 &
    reducedPartials_reducedPartials_carry_298; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_250 = reducedPartials_reducedPartials_sum_249 ^
    reducedPartials_reducedPartials_carry_297 ^ reducedPartials_reducedPartials_36_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_305 = reducedPartials_reducedPartials_sum_249 &
    reducedPartials_reducedPartials_carry_297 | reducedPartials_reducedPartials_carry_297 &
    reducedPartials_reducedPartials_36_0_1 | reducedPartials_reducedPartials_sum_249 &
    reducedPartials_reducedPartials_36_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_251 = reducedPartials_reducedPartials_sum_250 ^ partials_36_9 ^
    partials_36_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_306 = reducedPartials_reducedPartials_sum_250 & partials_36_9 |
    partials_36_9 & partials_36_10 | reducedPartials_reducedPartials_sum_250 & partials_36_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_252 = reducedPartials_reducedPartials_sum_251 ^ partials_36_11 ^
    partials_36_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_307 = reducedPartials_reducedPartials_sum_251 & partials_36_11 |
    partials_36_11 & partials_36_12 | reducedPartials_reducedPartials_sum_251 & partials_36_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_36_0_2 = reducedPartials_reducedPartials_sum_252 ^ partials_36_13 ^
    partials_36_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_308 = reducedPartials_reducedPartials_sum_252 & partials_36_13 |
    partials_36_13 & partials_36_14 | reducedPartials_reducedPartials_sum_252 & partials_36_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_253 = reducedPartials_reducedPartials_carry_308 ^
    reducedPartials_reducedPartials_carry_307 ^ reducedPartials_reducedPartials_carry_306; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_309 = reducedPartials_reducedPartials_carry_308 &
    reducedPartials_reducedPartials_carry_307 | reducedPartials_reducedPartials_carry_307 &
    reducedPartials_reducedPartials_carry_306 | reducedPartials_reducedPartials_carry_308 &
    reducedPartials_reducedPartials_carry_306; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_254 = reducedPartials_reducedPartials_sum_253 ^
    reducedPartials_reducedPartials_carry_305 ^ reducedPartials_reducedPartials_carry_304; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_310 = reducedPartials_reducedPartials_sum_253 &
    reducedPartials_reducedPartials_carry_305 | reducedPartials_reducedPartials_carry_305 &
    reducedPartials_reducedPartials_carry_304 | reducedPartials_reducedPartials_sum_253 &
    reducedPartials_reducedPartials_carry_304; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_255 = reducedPartials_reducedPartials_sum_254 ^
    reducedPartials_reducedPartials_carry_303 ^ reducedPartials_reducedPartials_37_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_311 = reducedPartials_reducedPartials_sum_254 &
    reducedPartials_reducedPartials_carry_303 | reducedPartials_reducedPartials_carry_303 &
    reducedPartials_reducedPartials_37_0 | reducedPartials_reducedPartials_sum_254 &
    reducedPartials_reducedPartials_37_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_256 = reducedPartials_reducedPartials_sum_255 ^ partials_37_8 ^
    partials_37_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_312 = reducedPartials_reducedPartials_sum_255 & partials_37_8 |
    partials_37_8 & partials_37_9 | reducedPartials_reducedPartials_sum_255 & partials_37_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_257 = reducedPartials_reducedPartials_sum_256 ^ partials_37_10 ^
    partials_37_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_313 = reducedPartials_reducedPartials_sum_256 & partials_37_10 |
    partials_37_10 & partials_37_11 | reducedPartials_reducedPartials_sum_256 & partials_37_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_37_0_1 = reducedPartials_reducedPartials_sum_257 ^ partials_37_12 ^
    partials_37_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_314 = reducedPartials_reducedPartials_sum_257 & partials_37_12 |
    partials_37_12 & partials_37_13 | reducedPartials_reducedPartials_sum_257 & partials_37_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_258 = reducedPartials_reducedPartials_carry_314 ^
    reducedPartials_reducedPartials_carry_313 ^ reducedPartials_reducedPartials_carry_312; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_315 = reducedPartials_reducedPartials_carry_314 &
    reducedPartials_reducedPartials_carry_313 | reducedPartials_reducedPartials_carry_313 &
    reducedPartials_reducedPartials_carry_312 | reducedPartials_reducedPartials_carry_314 &
    reducedPartials_reducedPartials_carry_312; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_259 = reducedPartials_reducedPartials_sum_258 ^
    reducedPartials_reducedPartials_carry_311 ^ reducedPartials_reducedPartials_carry_310; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_316 = reducedPartials_reducedPartials_sum_258 &
    reducedPartials_reducedPartials_carry_311 | reducedPartials_reducedPartials_carry_311 &
    reducedPartials_reducedPartials_carry_310 | reducedPartials_reducedPartials_sum_258 &
    reducedPartials_reducedPartials_carry_310; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_260 = reducedPartials_reducedPartials_sum_259 ^
    reducedPartials_reducedPartials_carry_309 ^ reducedPartials_reducedPartials_38_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_317 = reducedPartials_reducedPartials_sum_259 &
    reducedPartials_reducedPartials_carry_309 | reducedPartials_reducedPartials_carry_309 &
    reducedPartials_reducedPartials_38_0 | reducedPartials_reducedPartials_sum_259 &
    reducedPartials_reducedPartials_38_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_261 = reducedPartials_reducedPartials_sum_260 ^ partials_38_7 ^
    partials_38_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_318 = reducedPartials_reducedPartials_sum_260 & partials_38_7 |
    partials_38_7 & partials_38_8 | reducedPartials_reducedPartials_sum_260 & partials_38_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_262 = reducedPartials_reducedPartials_sum_261 ^ partials_38_9 ^
    partials_38_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_319 = reducedPartials_reducedPartials_sum_261 & partials_38_9 |
    partials_38_9 & partials_38_10 | reducedPartials_reducedPartials_sum_261 & partials_38_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_38_0_1 = reducedPartials_reducedPartials_sum_262 ^ partials_38_11 ^
    partials_38_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_320 = reducedPartials_reducedPartials_sum_262 & partials_38_11 |
    partials_38_11 & partials_38_12 | reducedPartials_reducedPartials_sum_262 & partials_38_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_263 = reducedPartials_reducedPartials_carry_320 ^
    reducedPartials_reducedPartials_carry_319 ^ reducedPartials_reducedPartials_carry_318; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_321 = reducedPartials_reducedPartials_carry_320 &
    reducedPartials_reducedPartials_carry_319 | reducedPartials_reducedPartials_carry_319 &
    reducedPartials_reducedPartials_carry_318 | reducedPartials_reducedPartials_carry_320 &
    reducedPartials_reducedPartials_carry_318; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_264 = reducedPartials_reducedPartials_sum_263 ^
    reducedPartials_reducedPartials_carry_317 ^ reducedPartials_reducedPartials_carry_316; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_322 = reducedPartials_reducedPartials_sum_263 &
    reducedPartials_reducedPartials_carry_317 | reducedPartials_reducedPartials_carry_317 &
    reducedPartials_reducedPartials_carry_316 | reducedPartials_reducedPartials_sum_263 &
    reducedPartials_reducedPartials_carry_316; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_265 = reducedPartials_reducedPartials_sum_264 ^
    reducedPartials_reducedPartials_carry_315 ^ reducedPartials_reducedPartials_39_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_323 = reducedPartials_reducedPartials_sum_264 &
    reducedPartials_reducedPartials_carry_315 | reducedPartials_reducedPartials_carry_315 &
    reducedPartials_reducedPartials_39_0 | reducedPartials_reducedPartials_sum_264 &
    reducedPartials_reducedPartials_39_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_266 = reducedPartials_reducedPartials_sum_265 ^ partials_39_6 ^
    partials_39_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_324 = reducedPartials_reducedPartials_sum_265 & partials_39_6 |
    partials_39_6 & partials_39_7 | reducedPartials_reducedPartials_sum_265 & partials_39_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_267 = reducedPartials_reducedPartials_sum_266 ^ partials_39_8 ^
    partials_39_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_325 = reducedPartials_reducedPartials_sum_266 & partials_39_8 |
    partials_39_8 & partials_39_9 | reducedPartials_reducedPartials_sum_266 & partials_39_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_39_0_1 = reducedPartials_reducedPartials_sum_267 ^ partials_39_10 ^
    partials_39_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_326 = reducedPartials_reducedPartials_sum_267 & partials_39_10 |
    partials_39_10 & partials_39_11 | reducedPartials_reducedPartials_sum_267 & partials_39_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_268 = reducedPartials_reducedPartials_carry_326 ^
    reducedPartials_reducedPartials_carry_325 ^ reducedPartials_reducedPartials_carry_324; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_327 = reducedPartials_reducedPartials_carry_326 &
    reducedPartials_reducedPartials_carry_325 | reducedPartials_reducedPartials_carry_325 &
    reducedPartials_reducedPartials_carry_324 | reducedPartials_reducedPartials_carry_326 &
    reducedPartials_reducedPartials_carry_324; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_269 = reducedPartials_reducedPartials_sum_268 ^
    reducedPartials_reducedPartials_carry_323 ^ reducedPartials_reducedPartials_carry_322; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_328 = reducedPartials_reducedPartials_sum_268 &
    reducedPartials_reducedPartials_carry_323 | reducedPartials_reducedPartials_carry_323 &
    reducedPartials_reducedPartials_carry_322 | reducedPartials_reducedPartials_sum_268 &
    reducedPartials_reducedPartials_carry_322; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_270 = reducedPartials_reducedPartials_sum_269 ^
    reducedPartials_reducedPartials_carry_321 ^ reducedPartials_reducedPartials_40_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_329 = reducedPartials_reducedPartials_sum_269 &
    reducedPartials_reducedPartials_carry_321 | reducedPartials_reducedPartials_carry_321 &
    reducedPartials_reducedPartials_40_0 | reducedPartials_reducedPartials_sum_269 &
    reducedPartials_reducedPartials_40_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_271 = reducedPartials_reducedPartials_sum_270 ^ partials_40_5 ^
    partials_40_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_330 = reducedPartials_reducedPartials_sum_270 & partials_40_5 |
    partials_40_5 & partials_40_6 | reducedPartials_reducedPartials_sum_270 & partials_40_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_272 = reducedPartials_reducedPartials_sum_271 ^ partials_40_7 ^
    partials_40_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_331 = reducedPartials_reducedPartials_sum_271 & partials_40_7 |
    partials_40_7 & partials_40_8 | reducedPartials_reducedPartials_sum_271 & partials_40_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_40_0_1 = reducedPartials_reducedPartials_sum_272 ^ partials_40_9 ^
    partials_40_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_332 = reducedPartials_reducedPartials_sum_272 & partials_40_9 |
    partials_40_9 & partials_40_10 | reducedPartials_reducedPartials_sum_272 & partials_40_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_273 = reducedPartials_reducedPartials_carry_332 ^
    reducedPartials_reducedPartials_carry_331 ^ reducedPartials_reducedPartials_carry_330; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_333 = reducedPartials_reducedPartials_carry_332 &
    reducedPartials_reducedPartials_carry_331 | reducedPartials_reducedPartials_carry_331 &
    reducedPartials_reducedPartials_carry_330 | reducedPartials_reducedPartials_carry_332 &
    reducedPartials_reducedPartials_carry_330; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_274 = reducedPartials_reducedPartials_sum_273 ^
    reducedPartials_reducedPartials_carry_329 ^ reducedPartials_reducedPartials_carry_328; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_334 = reducedPartials_reducedPartials_sum_273 &
    reducedPartials_reducedPartials_carry_329 | reducedPartials_reducedPartials_carry_329 &
    reducedPartials_reducedPartials_carry_328 | reducedPartials_reducedPartials_sum_273 &
    reducedPartials_reducedPartials_carry_328; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_275 = reducedPartials_reducedPartials_sum_274 ^
    reducedPartials_reducedPartials_carry_327 ^ reducedPartials_reducedPartials_41_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_335 = reducedPartials_reducedPartials_sum_274 &
    reducedPartials_reducedPartials_carry_327 | reducedPartials_reducedPartials_carry_327 &
    reducedPartials_reducedPartials_41_0 | reducedPartials_reducedPartials_sum_274 &
    reducedPartials_reducedPartials_41_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_276 = reducedPartials_reducedPartials_sum_275 ^ partials_41_4 ^
    partials_41_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_336 = reducedPartials_reducedPartials_sum_275 & partials_41_4 |
    partials_41_4 & partials_41_5 | reducedPartials_reducedPartials_sum_275 & partials_41_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_277 = reducedPartials_reducedPartials_sum_276 ^ partials_41_6 ^
    partials_41_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_337 = reducedPartials_reducedPartials_sum_276 & partials_41_6 |
    partials_41_6 & partials_41_7 | reducedPartials_reducedPartials_sum_276 & partials_41_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_41_0_1 = reducedPartials_reducedPartials_sum_277 ^ partials_41_8 ^ partials_41_9
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_338 = reducedPartials_reducedPartials_sum_277 & partials_41_8 |
    partials_41_8 & partials_41_9 | reducedPartials_reducedPartials_sum_277 & partials_41_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_278 = reducedPartials_reducedPartials_carry_338 ^
    reducedPartials_reducedPartials_carry_337 ^ reducedPartials_reducedPartials_carry_336; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_339 = reducedPartials_reducedPartials_carry_338 &
    reducedPartials_reducedPartials_carry_337 | reducedPartials_reducedPartials_carry_337 &
    reducedPartials_reducedPartials_carry_336 | reducedPartials_reducedPartials_carry_338 &
    reducedPartials_reducedPartials_carry_336; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_279 = reducedPartials_reducedPartials_sum_278 ^
    reducedPartials_reducedPartials_carry_335 ^ reducedPartials_reducedPartials_carry_334; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_340 = reducedPartials_reducedPartials_sum_278 &
    reducedPartials_reducedPartials_carry_335 | reducedPartials_reducedPartials_carry_335 &
    reducedPartials_reducedPartials_carry_334 | reducedPartials_reducedPartials_sum_278 &
    reducedPartials_reducedPartials_carry_334; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_280 = reducedPartials_reducedPartials_sum_279 ^
    reducedPartials_reducedPartials_carry_333 ^ reducedPartials_reducedPartials_42_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_341 = reducedPartials_reducedPartials_sum_279 &
    reducedPartials_reducedPartials_carry_333 | reducedPartials_reducedPartials_carry_333 &
    reducedPartials_reducedPartials_42_0 | reducedPartials_reducedPartials_sum_279 &
    reducedPartials_reducedPartials_42_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_281 = reducedPartials_reducedPartials_sum_280 ^ partials_42_3 ^
    partials_42_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_342 = reducedPartials_reducedPartials_sum_280 & partials_42_3 |
    partials_42_3 & partials_42_4 | reducedPartials_reducedPartials_sum_280 & partials_42_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_282 = reducedPartials_reducedPartials_sum_281 ^ partials_42_5 ^
    partials_42_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_343 = reducedPartials_reducedPartials_sum_281 & partials_42_5 |
    partials_42_5 & partials_42_6 | reducedPartials_reducedPartials_sum_281 & partials_42_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_42_0_1 = reducedPartials_reducedPartials_sum_282 ^ partials_42_7 ^ partials_42_8
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_344 = reducedPartials_reducedPartials_sum_282 & partials_42_7 |
    partials_42_7 & partials_42_8 | reducedPartials_reducedPartials_sum_282 & partials_42_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_283 = reducedPartials_reducedPartials_carry_344 ^
    reducedPartials_reducedPartials_carry_343 ^ reducedPartials_reducedPartials_carry_342; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_345 = reducedPartials_reducedPartials_carry_344 &
    reducedPartials_reducedPartials_carry_343 | reducedPartials_reducedPartials_carry_343 &
    reducedPartials_reducedPartials_carry_342 | reducedPartials_reducedPartials_carry_344 &
    reducedPartials_reducedPartials_carry_342; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_284 = reducedPartials_reducedPartials_sum_283 ^
    reducedPartials_reducedPartials_carry_341 ^ reducedPartials_reducedPartials_carry_340; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_346 = reducedPartials_reducedPartials_sum_283 &
    reducedPartials_reducedPartials_carry_341 | reducedPartials_reducedPartials_carry_341 &
    reducedPartials_reducedPartials_carry_340 | reducedPartials_reducedPartials_sum_283 &
    reducedPartials_reducedPartials_carry_340; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_285 = reducedPartials_reducedPartials_sum_284 ^
    reducedPartials_reducedPartials_carry_339 ^ reducedPartials_reducedPartials_43_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_347 = reducedPartials_reducedPartials_sum_284 &
    reducedPartials_reducedPartials_carry_339 | reducedPartials_reducedPartials_carry_339 &
    reducedPartials_reducedPartials_43_0 | reducedPartials_reducedPartials_sum_284 &
    reducedPartials_reducedPartials_43_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_286 = reducedPartials_reducedPartials_sum_285 ^ partials_43_2 ^
    partials_43_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_348 = reducedPartials_reducedPartials_sum_285 & partials_43_2 |
    partials_43_2 & partials_43_3 | reducedPartials_reducedPartials_sum_285 & partials_43_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_287 = reducedPartials_reducedPartials_sum_286 ^ partials_43_4 ^
    partials_43_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_349 = reducedPartials_reducedPartials_sum_286 & partials_43_4 |
    partials_43_4 & partials_43_5 | reducedPartials_reducedPartials_sum_286 & partials_43_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_43_0_1 = reducedPartials_reducedPartials_sum_287 ^ partials_43_6 ^ partials_43_7
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_350 = reducedPartials_reducedPartials_sum_287 & partials_43_6 |
    partials_43_6 & partials_43_7 | reducedPartials_reducedPartials_sum_287 & partials_43_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_288 = reducedPartials_reducedPartials_carry_350 ^
    reducedPartials_reducedPartials_carry_349 ^ reducedPartials_reducedPartials_carry_348; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_351 = reducedPartials_reducedPartials_carry_350 &
    reducedPartials_reducedPartials_carry_349 | reducedPartials_reducedPartials_carry_349 &
    reducedPartials_reducedPartials_carry_348 | reducedPartials_reducedPartials_carry_350 &
    reducedPartials_reducedPartials_carry_348; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_289 = reducedPartials_reducedPartials_sum_288 ^
    reducedPartials_reducedPartials_carry_347 ^ reducedPartials_reducedPartials_carry_346; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_352 = reducedPartials_reducedPartials_sum_288 &
    reducedPartials_reducedPartials_carry_347 | reducedPartials_reducedPartials_carry_347 &
    reducedPartials_reducedPartials_carry_346 | reducedPartials_reducedPartials_sum_288 &
    reducedPartials_reducedPartials_carry_346; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_290 = reducedPartials_reducedPartials_sum_289 ^
    reducedPartials_reducedPartials_carry_345 ^ reducedPartials_reducedPartials_44_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_353 = reducedPartials_reducedPartials_sum_289 &
    reducedPartials_reducedPartials_carry_345 | reducedPartials_reducedPartials_carry_345 &
    reducedPartials_reducedPartials_44_0 | reducedPartials_reducedPartials_sum_289 &
    reducedPartials_reducedPartials_44_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_291 = reducedPartials_reducedPartials_sum_290 ^ partials_44_1 ^
    partials_44_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_354 = reducedPartials_reducedPartials_sum_290 & partials_44_1 |
    partials_44_1 & partials_44_2 | reducedPartials_reducedPartials_sum_290 & partials_44_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_292 = reducedPartials_reducedPartials_sum_291 ^ partials_44_3 ^
    partials_44_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_355 = reducedPartials_reducedPartials_sum_291 & partials_44_3 |
    partials_44_3 & partials_44_4 | reducedPartials_reducedPartials_sum_291 & partials_44_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_44_0_1 = reducedPartials_reducedPartials_sum_292 ^ partials_44_5 ^ partials_44_6
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_356 = reducedPartials_reducedPartials_sum_292 & partials_44_5 |
    partials_44_5 & partials_44_6 | reducedPartials_reducedPartials_sum_292 & partials_44_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_293 = reducedPartials_reducedPartials_carry_356 ^
    reducedPartials_reducedPartials_carry_355 ^ reducedPartials_reducedPartials_carry_354; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_357 = reducedPartials_reducedPartials_carry_356 &
    reducedPartials_reducedPartials_carry_355 | reducedPartials_reducedPartials_carry_355 &
    reducedPartials_reducedPartials_carry_354 | reducedPartials_reducedPartials_carry_356 &
    reducedPartials_reducedPartials_carry_354; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_294 = reducedPartials_reducedPartials_sum_293 ^
    reducedPartials_reducedPartials_carry_353 ^ reducedPartials_reducedPartials_carry_352; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_358 = reducedPartials_reducedPartials_sum_293 &
    reducedPartials_reducedPartials_carry_353 | reducedPartials_reducedPartials_carry_353 &
    reducedPartials_reducedPartials_carry_352 | reducedPartials_reducedPartials_sum_293 &
    reducedPartials_reducedPartials_carry_352; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_295 = reducedPartials_reducedPartials_sum_294 ^
    reducedPartials_reducedPartials_carry_351 ^ reducedPartials_reducedPartials_45_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_359 = reducedPartials_reducedPartials_sum_294 &
    reducedPartials_reducedPartials_carry_351 | reducedPartials_reducedPartials_carry_351 &
    reducedPartials_reducedPartials_45_0 | reducedPartials_reducedPartials_sum_294 &
    reducedPartials_reducedPartials_45_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_296 = reducedPartials_reducedPartials_sum_295 ^ partials_45_0 ^
    partials_45_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_360 = reducedPartials_reducedPartials_sum_295 & partials_45_0 |
    partials_45_0 & partials_45_1 | reducedPartials_reducedPartials_sum_295 & partials_45_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_297 = reducedPartials_reducedPartials_sum_296 ^ partials_45_2 ^
    partials_45_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_361 = reducedPartials_reducedPartials_sum_296 & partials_45_2 |
    partials_45_2 & partials_45_3 | reducedPartials_reducedPartials_sum_296 & partials_45_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_45_0_1 = reducedPartials_reducedPartials_sum_297 ^ partials_45_4 ^ partials_45_5
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_362 = reducedPartials_reducedPartials_sum_297 & partials_45_4 |
    partials_45_4 & partials_45_5 | reducedPartials_reducedPartials_sum_297 & partials_45_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_298 = reducedPartials_reducedPartials_carry_362 ^
    reducedPartials_reducedPartials_carry_361 ^ reducedPartials_reducedPartials_carry_360; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_363 = reducedPartials_reducedPartials_carry_362 &
    reducedPartials_reducedPartials_carry_361 | reducedPartials_reducedPartials_carry_361 &
    reducedPartials_reducedPartials_carry_360 | reducedPartials_reducedPartials_carry_362 &
    reducedPartials_reducedPartials_carry_360; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_299 = reducedPartials_reducedPartials_sum_298 ^
    reducedPartials_reducedPartials_carry_359 ^ reducedPartials_reducedPartials_carry_358; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_364 = reducedPartials_reducedPartials_sum_298 &
    reducedPartials_reducedPartials_carry_359 | reducedPartials_reducedPartials_carry_359 &
    reducedPartials_reducedPartials_carry_358 | reducedPartials_reducedPartials_sum_298 &
    reducedPartials_reducedPartials_carry_358; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_300 = reducedPartials_reducedPartials_sum_299 ^
    reducedPartials_reducedPartials_carry_357 ^ partials_46_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_365 = reducedPartials_reducedPartials_sum_299 &
    reducedPartials_reducedPartials_carry_357 | reducedPartials_reducedPartials_carry_357 & partials_46_0 |
    reducedPartials_reducedPartials_sum_299 & partials_46_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_301 = reducedPartials_reducedPartials_sum_300 ^ partials_46_1 ^
    partials_46_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_366 = reducedPartials_reducedPartials_sum_300 & partials_46_1 |
    partials_46_1 & partials_46_2 | reducedPartials_reducedPartials_sum_300 & partials_46_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_46_0 = reducedPartials_reducedPartials_sum_301 ^ partials_46_3 ^ partials_46_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_367 = reducedPartials_reducedPartials_sum_301 & partials_46_3 |
    partials_46_3 & partials_46_4 | reducedPartials_reducedPartials_sum_301 & partials_46_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_302 = reducedPartials_reducedPartials_carry_367 ^
    reducedPartials_reducedPartials_carry_366 ^ reducedPartials_reducedPartials_carry_365; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_368 = reducedPartials_reducedPartials_carry_367 &
    reducedPartials_reducedPartials_carry_366 | reducedPartials_reducedPartials_carry_366 &
    reducedPartials_reducedPartials_carry_365 | reducedPartials_reducedPartials_carry_367 &
    reducedPartials_reducedPartials_carry_365; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_303 = reducedPartials_reducedPartials_sum_302 ^
    reducedPartials_reducedPartials_carry_364 ^ reducedPartials_reducedPartials_carry_363; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_369 = reducedPartials_reducedPartials_sum_302 &
    reducedPartials_reducedPartials_carry_364 | reducedPartials_reducedPartials_carry_364 &
    reducedPartials_reducedPartials_carry_363 | reducedPartials_reducedPartials_sum_302 &
    reducedPartials_reducedPartials_carry_363; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_304 = reducedPartials_reducedPartials_sum_303 ^ partials_47_0 ^
    partials_47_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_370 = reducedPartials_reducedPartials_sum_303 & partials_47_0 |
    partials_47_0 & partials_47_1 | reducedPartials_reducedPartials_sum_303 & partials_47_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_47_0 = reducedPartials_reducedPartials_sum_304 ^ partials_47_2 ^ partials_47_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_371 = reducedPartials_reducedPartials_sum_304 & partials_47_2 |
    partials_47_2 & partials_47_3 | reducedPartials_reducedPartials_sum_304 & partials_47_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_305 = reducedPartials_reducedPartials_carry_371 ^
    reducedPartials_reducedPartials_carry_370 ^ reducedPartials_reducedPartials_carry_369; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_372 = reducedPartials_reducedPartials_carry_371 &
    reducedPartials_reducedPartials_carry_370 | reducedPartials_reducedPartials_carry_370 &
    reducedPartials_reducedPartials_carry_369 | reducedPartials_reducedPartials_carry_371 &
    reducedPartials_reducedPartials_carry_369; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_306 = reducedPartials_reducedPartials_sum_305 ^
    reducedPartials_reducedPartials_carry_368 ^ partials_48_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_373 = reducedPartials_reducedPartials_sum_305 &
    reducedPartials_reducedPartials_carry_368 | reducedPartials_reducedPartials_carry_368 & partials_48_0 |
    reducedPartials_reducedPartials_sum_305 & partials_48_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_48_0 = reducedPartials_reducedPartials_sum_306 ^ partials_48_1 ^ partials_48_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_374 = reducedPartials_reducedPartials_sum_306 & partials_48_1 |
    partials_48_1 & partials_48_2 | reducedPartials_reducedPartials_sum_306 & partials_48_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_307 = reducedPartials_reducedPartials_carry_374 ^
    reducedPartials_reducedPartials_carry_373 ^ reducedPartials_reducedPartials_carry_372; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_375 = reducedPartials_reducedPartials_carry_374 &
    reducedPartials_reducedPartials_carry_373 | reducedPartials_reducedPartials_carry_373 &
    reducedPartials_reducedPartials_carry_372 | reducedPartials_reducedPartials_carry_374 &
    reducedPartials_reducedPartials_carry_372; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_49_0 = reducedPartials_reducedPartials_sum_307 ^ partials_49_0 ^ partials_49_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_376 = reducedPartials_reducedPartials_sum_307 & partials_49_0 |
    partials_49_0 & partials_49_1 | reducedPartials_reducedPartials_sum_307 & partials_49_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_50_0 = reducedPartials_reducedPartials_carry_376 ^
    reducedPartials_reducedPartials_carry_375 ^ partials_50_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_51_0 = reducedPartials_reducedPartials_carry_376 &
    reducedPartials_reducedPartials_carry_375 | reducedPartials_reducedPartials_carry_375 & partials_50_0 |
    reducedPartials_reducedPartials_carry_376 & partials_50_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_9_0 = partials_9_0 ^ partials_9_1; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_377 = partials_9_0 & partials_9_1; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_308 = reducedPartials_reducedPartials_carry_377 ^ partials_10_0 ^
    partials_10_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_378 = reducedPartials_reducedPartials_carry_377 & partials_10_0 |
    partials_10_0 & partials_10_1 | reducedPartials_reducedPartials_carry_377 & partials_10_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_10_0 = reducedPartials_reducedPartials_sum_308 ^ partials_10_2; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_379 = reducedPartials_reducedPartials_sum_308 & partials_10_2; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_309 = reducedPartials_reducedPartials_carry_379 ^
    reducedPartials_reducedPartials_carry_378 ^ partials_11_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_380 = reducedPartials_reducedPartials_carry_379 &
    reducedPartials_reducedPartials_carry_378 | reducedPartials_reducedPartials_carry_378 & partials_11_0 |
    reducedPartials_reducedPartials_carry_379 & partials_11_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_310 = reducedPartials_reducedPartials_sum_309 ^ partials_11_1 ^
    partials_11_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_381 = reducedPartials_reducedPartials_sum_309 & partials_11_1 |
    partials_11_1 & partials_11_2 | reducedPartials_reducedPartials_sum_309 & partials_11_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_11_0 = reducedPartials_reducedPartials_sum_310 ^ partials_11_3; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_382 = reducedPartials_reducedPartials_sum_310 & partials_11_3; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_311 = reducedPartials_reducedPartials_carry_382 ^
    reducedPartials_reducedPartials_carry_381 ^ reducedPartials_reducedPartials_carry_380; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_383 = reducedPartials_reducedPartials_carry_382 &
    reducedPartials_reducedPartials_carry_381 | reducedPartials_reducedPartials_carry_381 &
    reducedPartials_reducedPartials_carry_380 | reducedPartials_reducedPartials_carry_382 &
    reducedPartials_reducedPartials_carry_380; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_312 = reducedPartials_reducedPartials_sum_311 ^ partials_12_0 ^
    partials_12_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_384 = reducedPartials_reducedPartials_sum_311 & partials_12_0 |
    partials_12_0 & partials_12_1 | reducedPartials_reducedPartials_sum_311 & partials_12_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_313 = reducedPartials_reducedPartials_sum_312 ^ partials_12_2 ^
    partials_12_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_385 = reducedPartials_reducedPartials_sum_312 & partials_12_2 |
    partials_12_2 & partials_12_3 | reducedPartials_reducedPartials_sum_312 & partials_12_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_12_0 = reducedPartials_reducedPartials_sum_313 ^ partials_12_4; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_386 = reducedPartials_reducedPartials_sum_313 & partials_12_4; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_314 = reducedPartials_reducedPartials_carry_386 ^
    reducedPartials_reducedPartials_carry_385 ^ reducedPartials_reducedPartials_carry_384; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_387 = reducedPartials_reducedPartials_carry_386 &
    reducedPartials_reducedPartials_carry_385 | reducedPartials_reducedPartials_carry_385 &
    reducedPartials_reducedPartials_carry_384 | reducedPartials_reducedPartials_carry_386 &
    reducedPartials_reducedPartials_carry_384; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_315 = reducedPartials_reducedPartials_sum_314 ^
    reducedPartials_reducedPartials_carry_383 ^ reducedPartials_reducedPartials_13_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_388 = reducedPartials_reducedPartials_sum_314 &
    reducedPartials_reducedPartials_carry_383 | reducedPartials_reducedPartials_carry_383 &
    reducedPartials_reducedPartials_13_0 | reducedPartials_reducedPartials_sum_314 &
    reducedPartials_reducedPartials_13_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_316 = reducedPartials_reducedPartials_sum_315 ^ partials_13_2 ^
    partials_13_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_389 = reducedPartials_reducedPartials_sum_315 & partials_13_2 |
    partials_13_2 & partials_13_3 | reducedPartials_reducedPartials_sum_315 & partials_13_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_13_0_1 = reducedPartials_reducedPartials_sum_316 ^ partials_13_4 ^ partials_13_5
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_390 = reducedPartials_reducedPartials_sum_316 & partials_13_4 |
    partials_13_4 & partials_13_5 | reducedPartials_reducedPartials_sum_316 & partials_13_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_317 = reducedPartials_reducedPartials_carry_390 ^
    reducedPartials_reducedPartials_carry_389 ^ reducedPartials_reducedPartials_carry_388; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_391 = reducedPartials_reducedPartials_carry_390 &
    reducedPartials_reducedPartials_carry_389 | reducedPartials_reducedPartials_carry_389 &
    reducedPartials_reducedPartials_carry_388 | reducedPartials_reducedPartials_carry_390 &
    reducedPartials_reducedPartials_carry_388; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_318 = reducedPartials_reducedPartials_sum_317 ^
    reducedPartials_reducedPartials_carry_387 ^ reducedPartials_reducedPartials_14_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_392 = reducedPartials_reducedPartials_sum_317 &
    reducedPartials_reducedPartials_carry_387 | reducedPartials_reducedPartials_carry_387 &
    reducedPartials_reducedPartials_14_0 | reducedPartials_reducedPartials_sum_317 &
    reducedPartials_reducedPartials_14_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_319 = reducedPartials_reducedPartials_sum_318 ^ partials_14_3 ^
    partials_14_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_393 = reducedPartials_reducedPartials_sum_318 & partials_14_3 |
    partials_14_3 & partials_14_4 | reducedPartials_reducedPartials_sum_318 & partials_14_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_14_0_1 = reducedPartials_reducedPartials_sum_319 ^ partials_14_5 ^ partials_14_6
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_394 = reducedPartials_reducedPartials_sum_319 & partials_14_5 |
    partials_14_5 & partials_14_6 | reducedPartials_reducedPartials_sum_319 & partials_14_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_320 = reducedPartials_reducedPartials_carry_394 ^
    reducedPartials_reducedPartials_carry_393 ^ reducedPartials_reducedPartials_carry_392; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_395 = reducedPartials_reducedPartials_carry_394 &
    reducedPartials_reducedPartials_carry_393 | reducedPartials_reducedPartials_carry_393 &
    reducedPartials_reducedPartials_carry_392 | reducedPartials_reducedPartials_carry_394 &
    reducedPartials_reducedPartials_carry_392; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_321 = reducedPartials_reducedPartials_sum_320 ^
    reducedPartials_reducedPartials_carry_391 ^ reducedPartials_reducedPartials_15_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_396 = reducedPartials_reducedPartials_sum_320 &
    reducedPartials_reducedPartials_carry_391 | reducedPartials_reducedPartials_carry_391 &
    reducedPartials_reducedPartials_15_0 | reducedPartials_reducedPartials_sum_320 &
    reducedPartials_reducedPartials_15_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_322 = reducedPartials_reducedPartials_sum_321 ^ partials_15_4 ^
    partials_15_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_397 = reducedPartials_reducedPartials_sum_321 & partials_15_4 |
    partials_15_4 & partials_15_5 | reducedPartials_reducedPartials_sum_321 & partials_15_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_15_0_1 = reducedPartials_reducedPartials_sum_322 ^ partials_15_6 ^ partials_15_7
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_398 = reducedPartials_reducedPartials_sum_322 & partials_15_6 |
    partials_15_6 & partials_15_7 | reducedPartials_reducedPartials_sum_322 & partials_15_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_323 = reducedPartials_reducedPartials_carry_398 ^
    reducedPartials_reducedPartials_carry_397 ^ reducedPartials_reducedPartials_carry_396; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_399 = reducedPartials_reducedPartials_carry_398 &
    reducedPartials_reducedPartials_carry_397 | reducedPartials_reducedPartials_carry_397 &
    reducedPartials_reducedPartials_carry_396 | reducedPartials_reducedPartials_carry_398 &
    reducedPartials_reducedPartials_carry_396; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_324 = reducedPartials_reducedPartials_sum_323 ^
    reducedPartials_reducedPartials_carry_395 ^ reducedPartials_reducedPartials_16_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_400 = reducedPartials_reducedPartials_sum_323 &
    reducedPartials_reducedPartials_carry_395 | reducedPartials_reducedPartials_carry_395 &
    reducedPartials_reducedPartials_16_0 | reducedPartials_reducedPartials_sum_323 &
    reducedPartials_reducedPartials_16_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_325 = reducedPartials_reducedPartials_sum_324 ^ partials_16_5 ^
    partials_16_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_401 = reducedPartials_reducedPartials_sum_324 & partials_16_5 |
    partials_16_5 & partials_16_6 | reducedPartials_reducedPartials_sum_324 & partials_16_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_16_0_1 = reducedPartials_reducedPartials_sum_325 ^ partials_16_7 ^ partials_16_8
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_402 = reducedPartials_reducedPartials_sum_325 & partials_16_7 |
    partials_16_7 & partials_16_8 | reducedPartials_reducedPartials_sum_325 & partials_16_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_326 = reducedPartials_reducedPartials_carry_402 ^
    reducedPartials_reducedPartials_carry_401 ^ reducedPartials_reducedPartials_carry_400; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_403 = reducedPartials_reducedPartials_carry_402 &
    reducedPartials_reducedPartials_carry_401 | reducedPartials_reducedPartials_carry_401 &
    reducedPartials_reducedPartials_carry_400 | reducedPartials_reducedPartials_carry_402 &
    reducedPartials_reducedPartials_carry_400; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_327 = reducedPartials_reducedPartials_sum_326 ^
    reducedPartials_reducedPartials_carry_399 ^ reducedPartials_reducedPartials_17_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_404 = reducedPartials_reducedPartials_sum_326 &
    reducedPartials_reducedPartials_carry_399 | reducedPartials_reducedPartials_carry_399 &
    reducedPartials_reducedPartials_17_0 | reducedPartials_reducedPartials_sum_326 &
    reducedPartials_reducedPartials_17_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_328 = reducedPartials_reducedPartials_sum_327 ^ partials_17_6 ^
    partials_17_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_405 = reducedPartials_reducedPartials_sum_327 & partials_17_6 |
    partials_17_6 & partials_17_7 | reducedPartials_reducedPartials_sum_327 & partials_17_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_17_0_1 = reducedPartials_reducedPartials_sum_328 ^ partials_17_8 ^ partials_17_9
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_406 = reducedPartials_reducedPartials_sum_328 & partials_17_8 |
    partials_17_8 & partials_17_9 | reducedPartials_reducedPartials_sum_328 & partials_17_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_329 = reducedPartials_reducedPartials_carry_406 ^
    reducedPartials_reducedPartials_carry_405 ^ reducedPartials_reducedPartials_carry_404; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_407 = reducedPartials_reducedPartials_carry_406 &
    reducedPartials_reducedPartials_carry_405 | reducedPartials_reducedPartials_carry_405 &
    reducedPartials_reducedPartials_carry_404 | reducedPartials_reducedPartials_carry_406 &
    reducedPartials_reducedPartials_carry_404; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_330 = reducedPartials_reducedPartials_sum_329 ^
    reducedPartials_reducedPartials_carry_403 ^ reducedPartials_reducedPartials_18_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_408 = reducedPartials_reducedPartials_sum_329 &
    reducedPartials_reducedPartials_carry_403 | reducedPartials_reducedPartials_carry_403 &
    reducedPartials_reducedPartials_18_0 | reducedPartials_reducedPartials_sum_329 &
    reducedPartials_reducedPartials_18_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_331 = reducedPartials_reducedPartials_sum_330 ^ partials_18_7 ^
    partials_18_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_409 = reducedPartials_reducedPartials_sum_330 & partials_18_7 |
    partials_18_7 & partials_18_8 | reducedPartials_reducedPartials_sum_330 & partials_18_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_18_0_1 = reducedPartials_reducedPartials_sum_331 ^ partials_18_9 ^
    partials_18_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_410 = reducedPartials_reducedPartials_sum_331 & partials_18_9 |
    partials_18_9 & partials_18_10 | reducedPartials_reducedPartials_sum_331 & partials_18_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_332 = reducedPartials_reducedPartials_carry_410 ^
    reducedPartials_reducedPartials_carry_409 ^ reducedPartials_reducedPartials_carry_408; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_411 = reducedPartials_reducedPartials_carry_410 &
    reducedPartials_reducedPartials_carry_409 | reducedPartials_reducedPartials_carry_409 &
    reducedPartials_reducedPartials_carry_408 | reducedPartials_reducedPartials_carry_410 &
    reducedPartials_reducedPartials_carry_408; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_333 = reducedPartials_reducedPartials_sum_332 ^
    reducedPartials_reducedPartials_carry_407 ^ reducedPartials_reducedPartials_19_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_412 = reducedPartials_reducedPartials_sum_332 &
    reducedPartials_reducedPartials_carry_407 | reducedPartials_reducedPartials_carry_407 &
    reducedPartials_reducedPartials_19_0_1 | reducedPartials_reducedPartials_sum_332 &
    reducedPartials_reducedPartials_19_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_334 = reducedPartials_reducedPartials_sum_333 ^ partials_19_8 ^
    partials_19_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_413 = reducedPartials_reducedPartials_sum_333 & partials_19_8 |
    partials_19_8 & partials_19_9 | reducedPartials_reducedPartials_sum_333 & partials_19_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_19_0_2 = reducedPartials_reducedPartials_sum_334 ^ partials_19_10 ^
    partials_19_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_414 = reducedPartials_reducedPartials_sum_334 & partials_19_10 |
    partials_19_10 & partials_19_11 | reducedPartials_reducedPartials_sum_334 & partials_19_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_335 = reducedPartials_reducedPartials_carry_414 ^
    reducedPartials_reducedPartials_carry_413 ^ reducedPartials_reducedPartials_carry_412; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_415 = reducedPartials_reducedPartials_carry_414 &
    reducedPartials_reducedPartials_carry_413 | reducedPartials_reducedPartials_carry_413 &
    reducedPartials_reducedPartials_carry_412 | reducedPartials_reducedPartials_carry_414 &
    reducedPartials_reducedPartials_carry_412; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_336 = reducedPartials_reducedPartials_sum_335 ^
    reducedPartials_reducedPartials_carry_411 ^ reducedPartials_reducedPartials_20_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_416 = reducedPartials_reducedPartials_sum_335 &
    reducedPartials_reducedPartials_carry_411 | reducedPartials_reducedPartials_carry_411 &
    reducedPartials_reducedPartials_20_0_1 | reducedPartials_reducedPartials_sum_335 &
    reducedPartials_reducedPartials_20_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_337 = reducedPartials_reducedPartials_sum_336 ^ partials_20_9 ^
    partials_20_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_417 = reducedPartials_reducedPartials_sum_336 & partials_20_9 |
    partials_20_9 & partials_20_10 | reducedPartials_reducedPartials_sum_336 & partials_20_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_20_0_2 = reducedPartials_reducedPartials_sum_337 ^ partials_20_11 ^
    partials_20_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_418 = reducedPartials_reducedPartials_sum_337 & partials_20_11 |
    partials_20_11 & partials_20_12 | reducedPartials_reducedPartials_sum_337 & partials_20_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_338 = reducedPartials_reducedPartials_carry_418 ^
    reducedPartials_reducedPartials_carry_417 ^ reducedPartials_reducedPartials_carry_416; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_419 = reducedPartials_reducedPartials_carry_418 &
    reducedPartials_reducedPartials_carry_417 | reducedPartials_reducedPartials_carry_417 &
    reducedPartials_reducedPartials_carry_416 | reducedPartials_reducedPartials_carry_418 &
    reducedPartials_reducedPartials_carry_416; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_339 = reducedPartials_reducedPartials_sum_338 ^
    reducedPartials_reducedPartials_carry_415 ^ reducedPartials_reducedPartials_21_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_420 = reducedPartials_reducedPartials_sum_338 &
    reducedPartials_reducedPartials_carry_415 | reducedPartials_reducedPartials_carry_415 &
    reducedPartials_reducedPartials_21_0_1 | reducedPartials_reducedPartials_sum_338 &
    reducedPartials_reducedPartials_21_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_340 = reducedPartials_reducedPartials_sum_339 ^ partials_21_10 ^
    partials_21_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_421 = reducedPartials_reducedPartials_sum_339 & partials_21_10 |
    partials_21_10 & partials_21_11 | reducedPartials_reducedPartials_sum_339 & partials_21_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_21_0_2 = reducedPartials_reducedPartials_sum_340 ^ partials_21_12 ^
    partials_21_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_422 = reducedPartials_reducedPartials_sum_340 & partials_21_12 |
    partials_21_12 & partials_21_13 | reducedPartials_reducedPartials_sum_340 & partials_21_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_341 = reducedPartials_reducedPartials_carry_422 ^
    reducedPartials_reducedPartials_carry_421 ^ reducedPartials_reducedPartials_carry_420; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_423 = reducedPartials_reducedPartials_carry_422 &
    reducedPartials_reducedPartials_carry_421 | reducedPartials_reducedPartials_carry_421 &
    reducedPartials_reducedPartials_carry_420 | reducedPartials_reducedPartials_carry_422 &
    reducedPartials_reducedPartials_carry_420; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_342 = reducedPartials_reducedPartials_sum_341 ^
    reducedPartials_reducedPartials_carry_419 ^ reducedPartials_reducedPartials_22_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_424 = reducedPartials_reducedPartials_sum_341 &
    reducedPartials_reducedPartials_carry_419 | reducedPartials_reducedPartials_carry_419 &
    reducedPartials_reducedPartials_22_0_1 | reducedPartials_reducedPartials_sum_341 &
    reducedPartials_reducedPartials_22_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_343 = reducedPartials_reducedPartials_sum_342 ^ partials_22_11 ^
    partials_22_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_425 = reducedPartials_reducedPartials_sum_342 & partials_22_11 |
    partials_22_11 & partials_22_12 | reducedPartials_reducedPartials_sum_342 & partials_22_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_22_0_2 = reducedPartials_reducedPartials_sum_343 ^ partials_22_13 ^
    partials_22_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_426 = reducedPartials_reducedPartials_sum_343 & partials_22_13 |
    partials_22_13 & partials_22_14 | reducedPartials_reducedPartials_sum_343 & partials_22_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_344 = reducedPartials_reducedPartials_carry_426 ^
    reducedPartials_reducedPartials_carry_425 ^ reducedPartials_reducedPartials_carry_424; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_427 = reducedPartials_reducedPartials_carry_426 &
    reducedPartials_reducedPartials_carry_425 | reducedPartials_reducedPartials_carry_425 &
    reducedPartials_reducedPartials_carry_424 | reducedPartials_reducedPartials_carry_426 &
    reducedPartials_reducedPartials_carry_424; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_345 = reducedPartials_reducedPartials_sum_344 ^
    reducedPartials_reducedPartials_carry_423 ^ reducedPartials_reducedPartials_23_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_428 = reducedPartials_reducedPartials_sum_344 &
    reducedPartials_reducedPartials_carry_423 | reducedPartials_reducedPartials_carry_423 &
    reducedPartials_reducedPartials_23_0_1 | reducedPartials_reducedPartials_sum_344 &
    reducedPartials_reducedPartials_23_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_346 = reducedPartials_reducedPartials_sum_345 ^ partials_23_12 ^
    partials_23_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_429 = reducedPartials_reducedPartials_sum_345 & partials_23_12 |
    partials_23_12 & partials_23_13 | reducedPartials_reducedPartials_sum_345 & partials_23_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_23_0_2 = reducedPartials_reducedPartials_sum_346 ^ partials_23_14 ^
    partials_23_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_430 = reducedPartials_reducedPartials_sum_346 & partials_23_14 |
    partials_23_14 & partials_23_15 | reducedPartials_reducedPartials_sum_346 & partials_23_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_347 = reducedPartials_reducedPartials_carry_430 ^
    reducedPartials_reducedPartials_carry_429 ^ reducedPartials_reducedPartials_carry_428; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_431 = reducedPartials_reducedPartials_carry_430 &
    reducedPartials_reducedPartials_carry_429 | reducedPartials_reducedPartials_carry_429 &
    reducedPartials_reducedPartials_carry_428 | reducedPartials_reducedPartials_carry_430 &
    reducedPartials_reducedPartials_carry_428; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_348 = reducedPartials_reducedPartials_sum_347 ^
    reducedPartials_reducedPartials_carry_427 ^ reducedPartials_reducedPartials_24_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_432 = reducedPartials_reducedPartials_sum_347 &
    reducedPartials_reducedPartials_carry_427 | reducedPartials_reducedPartials_carry_427 &
    reducedPartials_reducedPartials_24_0_1 | reducedPartials_reducedPartials_sum_347 &
    reducedPartials_reducedPartials_24_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_349 = reducedPartials_reducedPartials_sum_348 ^ partials_24_13 ^
    partials_24_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_433 = reducedPartials_reducedPartials_sum_348 & partials_24_13 |
    partials_24_13 & partials_24_14 | reducedPartials_reducedPartials_sum_348 & partials_24_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_24_0_2 = reducedPartials_reducedPartials_sum_349 ^ partials_24_15 ^
    partials_24_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_434 = reducedPartials_reducedPartials_sum_349 & partials_24_15 |
    partials_24_15 & partials_24_16 | reducedPartials_reducedPartials_sum_349 & partials_24_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_350 = reducedPartials_reducedPartials_carry_434 ^
    reducedPartials_reducedPartials_carry_433 ^ reducedPartials_reducedPartials_carry_432; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_435 = reducedPartials_reducedPartials_carry_434 &
    reducedPartials_reducedPartials_carry_433 | reducedPartials_reducedPartials_carry_433 &
    reducedPartials_reducedPartials_carry_432 | reducedPartials_reducedPartials_carry_434 &
    reducedPartials_reducedPartials_carry_432; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_351 = reducedPartials_reducedPartials_sum_350 ^
    reducedPartials_reducedPartials_carry_431 ^ reducedPartials_reducedPartials_25_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_436 = reducedPartials_reducedPartials_sum_350 &
    reducedPartials_reducedPartials_carry_431 | reducedPartials_reducedPartials_carry_431 &
    reducedPartials_reducedPartials_25_0_1 | reducedPartials_reducedPartials_sum_350 &
    reducedPartials_reducedPartials_25_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_352 = reducedPartials_reducedPartials_sum_351 ^ partials_25_14 ^
    partials_25_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_437 = reducedPartials_reducedPartials_sum_351 & partials_25_14 |
    partials_25_14 & partials_25_15 | reducedPartials_reducedPartials_sum_351 & partials_25_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_25_0_2 = reducedPartials_reducedPartials_sum_352 ^ partials_25_16 ^
    partials_25_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_438 = reducedPartials_reducedPartials_sum_352 & partials_25_16 |
    partials_25_16 & partials_25_17 | reducedPartials_reducedPartials_sum_352 & partials_25_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_353 = reducedPartials_reducedPartials_carry_438 ^
    reducedPartials_reducedPartials_carry_437 ^ reducedPartials_reducedPartials_carry_436; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_439 = reducedPartials_reducedPartials_carry_438 &
    reducedPartials_reducedPartials_carry_437 | reducedPartials_reducedPartials_carry_437 &
    reducedPartials_reducedPartials_carry_436 | reducedPartials_reducedPartials_carry_438 &
    reducedPartials_reducedPartials_carry_436; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_354 = reducedPartials_reducedPartials_sum_353 ^
    reducedPartials_reducedPartials_carry_435 ^ reducedPartials_reducedPartials_26_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_440 = reducedPartials_reducedPartials_sum_353 &
    reducedPartials_reducedPartials_carry_435 | reducedPartials_reducedPartials_carry_435 &
    reducedPartials_reducedPartials_26_0_1 | reducedPartials_reducedPartials_sum_353 &
    reducedPartials_reducedPartials_26_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_355 = reducedPartials_reducedPartials_sum_354 ^ partials_26_15 ^
    partials_26_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_441 = reducedPartials_reducedPartials_sum_354 & partials_26_15 |
    partials_26_15 & partials_26_16 | reducedPartials_reducedPartials_sum_354 & partials_26_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_26_0_2 = reducedPartials_reducedPartials_sum_355 ^ partials_26_17 ^
    partials_26_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_442 = reducedPartials_reducedPartials_sum_355 & partials_26_17 |
    partials_26_17 & partials_26_18 | reducedPartials_reducedPartials_sum_355 & partials_26_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_356 = reducedPartials_reducedPartials_carry_442 ^
    reducedPartials_reducedPartials_carry_441 ^ reducedPartials_reducedPartials_carry_440; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_443 = reducedPartials_reducedPartials_carry_442 &
    reducedPartials_reducedPartials_carry_441 | reducedPartials_reducedPartials_carry_441 &
    reducedPartials_reducedPartials_carry_440 | reducedPartials_reducedPartials_carry_442 &
    reducedPartials_reducedPartials_carry_440; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_357 = reducedPartials_reducedPartials_sum_356 ^
    reducedPartials_reducedPartials_carry_439 ^ reducedPartials_reducedPartials_27_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_444 = reducedPartials_reducedPartials_sum_356 &
    reducedPartials_reducedPartials_carry_439 | reducedPartials_reducedPartials_carry_439 &
    reducedPartials_reducedPartials_27_0_1 | reducedPartials_reducedPartials_sum_356 &
    reducedPartials_reducedPartials_27_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_358 = reducedPartials_reducedPartials_sum_357 ^ partials_27_16 ^
    partials_27_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_445 = reducedPartials_reducedPartials_sum_357 & partials_27_16 |
    partials_27_16 & partials_27_17 | reducedPartials_reducedPartials_sum_357 & partials_27_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_27_0_2 = reducedPartials_reducedPartials_sum_358 ^ partials_27_18 ^
    partials_27_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_446 = reducedPartials_reducedPartials_sum_358 & partials_27_18 |
    partials_27_18 & partials_27_19 | reducedPartials_reducedPartials_sum_358 & partials_27_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_359 = reducedPartials_reducedPartials_carry_446 ^
    reducedPartials_reducedPartials_carry_445 ^ reducedPartials_reducedPartials_carry_444; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_447 = reducedPartials_reducedPartials_carry_446 &
    reducedPartials_reducedPartials_carry_445 | reducedPartials_reducedPartials_carry_445 &
    reducedPartials_reducedPartials_carry_444 | reducedPartials_reducedPartials_carry_446 &
    reducedPartials_reducedPartials_carry_444; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_360 = reducedPartials_reducedPartials_sum_359 ^
    reducedPartials_reducedPartials_carry_443 ^ reducedPartials_reducedPartials_28_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_448 = reducedPartials_reducedPartials_sum_359 &
    reducedPartials_reducedPartials_carry_443 | reducedPartials_reducedPartials_carry_443 &
    reducedPartials_reducedPartials_28_0_2 | reducedPartials_reducedPartials_sum_359 &
    reducedPartials_reducedPartials_28_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_361 = reducedPartials_reducedPartials_sum_360 ^ partials_28_17 ^
    partials_28_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_449 = reducedPartials_reducedPartials_sum_360 & partials_28_17 |
    partials_28_17 & partials_28_18 | reducedPartials_reducedPartials_sum_360 & partials_28_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_28_0_3 = reducedPartials_reducedPartials_sum_361 ^ partials_28_19 ^
    partials_28_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_450 = reducedPartials_reducedPartials_sum_361 & partials_28_19 |
    partials_28_19 & partials_28_20 | reducedPartials_reducedPartials_sum_361 & partials_28_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_362 = reducedPartials_reducedPartials_carry_450 ^
    reducedPartials_reducedPartials_carry_449 ^ reducedPartials_reducedPartials_carry_448; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_451 = reducedPartials_reducedPartials_carry_450 &
    reducedPartials_reducedPartials_carry_449 | reducedPartials_reducedPartials_carry_449 &
    reducedPartials_reducedPartials_carry_448 | reducedPartials_reducedPartials_carry_450 &
    reducedPartials_reducedPartials_carry_448; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_363 = reducedPartials_reducedPartials_sum_362 ^
    reducedPartials_reducedPartials_carry_447 ^ reducedPartials_reducedPartials_29_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_452 = reducedPartials_reducedPartials_sum_362 &
    reducedPartials_reducedPartials_carry_447 | reducedPartials_reducedPartials_carry_447 &
    reducedPartials_reducedPartials_29_0_2 | reducedPartials_reducedPartials_sum_362 &
    reducedPartials_reducedPartials_29_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_364 = reducedPartials_reducedPartials_sum_363 ^ partials_29_18 ^
    partials_29_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_453 = reducedPartials_reducedPartials_sum_363 & partials_29_18 |
    partials_29_18 & partials_29_19 | reducedPartials_reducedPartials_sum_363 & partials_29_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_29_0_3 = reducedPartials_reducedPartials_sum_364 ^ partials_29_20 ^
    partials_29_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_454 = reducedPartials_reducedPartials_sum_364 & partials_29_20 |
    partials_29_20 & partials_29_21 | reducedPartials_reducedPartials_sum_364 & partials_29_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_365 = reducedPartials_reducedPartials_carry_454 ^
    reducedPartials_reducedPartials_carry_453 ^ reducedPartials_reducedPartials_carry_452; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_455 = reducedPartials_reducedPartials_carry_454 &
    reducedPartials_reducedPartials_carry_453 | reducedPartials_reducedPartials_carry_453 &
    reducedPartials_reducedPartials_carry_452 | reducedPartials_reducedPartials_carry_454 &
    reducedPartials_reducedPartials_carry_452; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_366 = reducedPartials_reducedPartials_sum_365 ^
    reducedPartials_reducedPartials_carry_451 ^ reducedPartials_reducedPartials_30_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_456 = reducedPartials_reducedPartials_sum_365 &
    reducedPartials_reducedPartials_carry_451 | reducedPartials_reducedPartials_carry_451 &
    reducedPartials_reducedPartials_30_0_2 | reducedPartials_reducedPartials_sum_365 &
    reducedPartials_reducedPartials_30_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_367 = reducedPartials_reducedPartials_sum_366 ^ partials_30_19 ^
    partials_30_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_457 = reducedPartials_reducedPartials_sum_366 & partials_30_19 |
    partials_30_19 & partials_30_20 | reducedPartials_reducedPartials_sum_366 & partials_30_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_30_0_3 = reducedPartials_reducedPartials_sum_367 ^ partials_30_21 ^
    partials_30_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_458 = reducedPartials_reducedPartials_sum_367 & partials_30_21 |
    partials_30_21 & partials_30_22 | reducedPartials_reducedPartials_sum_367 & partials_30_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_368 = reducedPartials_reducedPartials_carry_458 ^
    reducedPartials_reducedPartials_carry_457 ^ reducedPartials_reducedPartials_carry_456; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_459 = reducedPartials_reducedPartials_carry_458 &
    reducedPartials_reducedPartials_carry_457 | reducedPartials_reducedPartials_carry_457 &
    reducedPartials_reducedPartials_carry_456 | reducedPartials_reducedPartials_carry_458 &
    reducedPartials_reducedPartials_carry_456; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_369 = reducedPartials_reducedPartials_sum_368 ^
    reducedPartials_reducedPartials_carry_455 ^ reducedPartials_reducedPartials_31_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_460 = reducedPartials_reducedPartials_sum_368 &
    reducedPartials_reducedPartials_carry_455 | reducedPartials_reducedPartials_carry_455 &
    reducedPartials_reducedPartials_31_0_2 | reducedPartials_reducedPartials_sum_368 &
    reducedPartials_reducedPartials_31_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_370 = reducedPartials_reducedPartials_sum_369 ^ partials_31_20 ^
    partials_31_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_461 = reducedPartials_reducedPartials_sum_369 & partials_31_20 |
    partials_31_20 & partials_31_21 | reducedPartials_reducedPartials_sum_369 & partials_31_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_31_0_3 = reducedPartials_reducedPartials_sum_370 ^ partials_31_22 ^
    partials_31_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_462 = reducedPartials_reducedPartials_sum_370 & partials_31_22 |
    partials_31_22 & partials_31_23 | reducedPartials_reducedPartials_sum_370 & partials_31_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_371 = reducedPartials_reducedPartials_carry_462 ^
    reducedPartials_reducedPartials_carry_461 ^ reducedPartials_reducedPartials_carry_460; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_463 = reducedPartials_reducedPartials_carry_462 &
    reducedPartials_reducedPartials_carry_461 | reducedPartials_reducedPartials_carry_461 &
    reducedPartials_reducedPartials_carry_460 | reducedPartials_reducedPartials_carry_462 &
    reducedPartials_reducedPartials_carry_460; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_372 = reducedPartials_reducedPartials_sum_371 ^
    reducedPartials_reducedPartials_carry_459 ^ reducedPartials_reducedPartials_32_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_464 = reducedPartials_reducedPartials_sum_371 &
    reducedPartials_reducedPartials_carry_459 | reducedPartials_reducedPartials_carry_459 &
    reducedPartials_reducedPartials_32_0_2 | reducedPartials_reducedPartials_sum_371 &
    reducedPartials_reducedPartials_32_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_373 = reducedPartials_reducedPartials_sum_372 ^ partials_32_19 ^
    partials_32_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_465 = reducedPartials_reducedPartials_sum_372 & partials_32_19 |
    partials_32_19 & partials_32_20 | reducedPartials_reducedPartials_sum_372 & partials_32_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_32_0_3 = reducedPartials_reducedPartials_sum_373 ^ partials_32_21 ^
    partials_32_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_466 = reducedPartials_reducedPartials_sum_373 & partials_32_21 |
    partials_32_21 & partials_32_22 | reducedPartials_reducedPartials_sum_373 & partials_32_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_374 = reducedPartials_reducedPartials_carry_466 ^
    reducedPartials_reducedPartials_carry_465 ^ reducedPartials_reducedPartials_carry_464; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_467 = reducedPartials_reducedPartials_carry_466 &
    reducedPartials_reducedPartials_carry_465 | reducedPartials_reducedPartials_carry_465 &
    reducedPartials_reducedPartials_carry_464 | reducedPartials_reducedPartials_carry_466 &
    reducedPartials_reducedPartials_carry_464; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_375 = reducedPartials_reducedPartials_sum_374 ^
    reducedPartials_reducedPartials_carry_463 ^ reducedPartials_reducedPartials_33_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_468 = reducedPartials_reducedPartials_sum_374 &
    reducedPartials_reducedPartials_carry_463 | reducedPartials_reducedPartials_carry_463 &
    reducedPartials_reducedPartials_33_0_2 | reducedPartials_reducedPartials_sum_374 &
    reducedPartials_reducedPartials_33_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_376 = reducedPartials_reducedPartials_sum_375 ^ partials_33_18 ^
    partials_33_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_469 = reducedPartials_reducedPartials_sum_375 & partials_33_18 |
    partials_33_18 & partials_33_19 | reducedPartials_reducedPartials_sum_375 & partials_33_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_33_0_3 = reducedPartials_reducedPartials_sum_376 ^ partials_33_20 ^
    partials_33_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_470 = reducedPartials_reducedPartials_sum_376 & partials_33_20 |
    partials_33_20 & partials_33_21 | reducedPartials_reducedPartials_sum_376 & partials_33_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_377 = reducedPartials_reducedPartials_carry_470 ^
    reducedPartials_reducedPartials_carry_469 ^ reducedPartials_reducedPartials_carry_468; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_471 = reducedPartials_reducedPartials_carry_470 &
    reducedPartials_reducedPartials_carry_469 | reducedPartials_reducedPartials_carry_469 &
    reducedPartials_reducedPartials_carry_468 | reducedPartials_reducedPartials_carry_470 &
    reducedPartials_reducedPartials_carry_468; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_378 = reducedPartials_reducedPartials_sum_377 ^
    reducedPartials_reducedPartials_carry_467 ^ reducedPartials_reducedPartials_34_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_472 = reducedPartials_reducedPartials_sum_377 &
    reducedPartials_reducedPartials_carry_467 | reducedPartials_reducedPartials_carry_467 &
    reducedPartials_reducedPartials_34_0_2 | reducedPartials_reducedPartials_sum_377 &
    reducedPartials_reducedPartials_34_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_379 = reducedPartials_reducedPartials_sum_378 ^ partials_34_17 ^
    partials_34_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_473 = reducedPartials_reducedPartials_sum_378 & partials_34_17 |
    partials_34_17 & partials_34_18 | reducedPartials_reducedPartials_sum_378 & partials_34_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_34_0_3 = reducedPartials_reducedPartials_sum_379 ^ partials_34_19 ^
    partials_34_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_474 = reducedPartials_reducedPartials_sum_379 & partials_34_19 |
    partials_34_19 & partials_34_20 | reducedPartials_reducedPartials_sum_379 & partials_34_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_380 = reducedPartials_reducedPartials_carry_474 ^
    reducedPartials_reducedPartials_carry_473 ^ reducedPartials_reducedPartials_carry_472; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_475 = reducedPartials_reducedPartials_carry_474 &
    reducedPartials_reducedPartials_carry_473 | reducedPartials_reducedPartials_carry_473 &
    reducedPartials_reducedPartials_carry_472 | reducedPartials_reducedPartials_carry_474 &
    reducedPartials_reducedPartials_carry_472; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_381 = reducedPartials_reducedPartials_sum_380 ^
    reducedPartials_reducedPartials_carry_471 ^ reducedPartials_reducedPartials_35_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_476 = reducedPartials_reducedPartials_sum_380 &
    reducedPartials_reducedPartials_carry_471 | reducedPartials_reducedPartials_carry_471 &
    reducedPartials_reducedPartials_35_0_2 | reducedPartials_reducedPartials_sum_380 &
    reducedPartials_reducedPartials_35_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_382 = reducedPartials_reducedPartials_sum_381 ^ partials_35_16 ^
    partials_35_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_477 = reducedPartials_reducedPartials_sum_381 & partials_35_16 |
    partials_35_16 & partials_35_17 | reducedPartials_reducedPartials_sum_381 & partials_35_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_35_0_3 = reducedPartials_reducedPartials_sum_382 ^ partials_35_18 ^
    partials_35_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_478 = reducedPartials_reducedPartials_sum_382 & partials_35_18 |
    partials_35_18 & partials_35_19 | reducedPartials_reducedPartials_sum_382 & partials_35_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_383 = reducedPartials_reducedPartials_carry_478 ^
    reducedPartials_reducedPartials_carry_477 ^ reducedPartials_reducedPartials_carry_476; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_479 = reducedPartials_reducedPartials_carry_478 &
    reducedPartials_reducedPartials_carry_477 | reducedPartials_reducedPartials_carry_477 &
    reducedPartials_reducedPartials_carry_476 | reducedPartials_reducedPartials_carry_478 &
    reducedPartials_reducedPartials_carry_476; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_384 = reducedPartials_reducedPartials_sum_383 ^
    reducedPartials_reducedPartials_carry_475 ^ reducedPartials_reducedPartials_36_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_480 = reducedPartials_reducedPartials_sum_383 &
    reducedPartials_reducedPartials_carry_475 | reducedPartials_reducedPartials_carry_475 &
    reducedPartials_reducedPartials_36_0_2 | reducedPartials_reducedPartials_sum_383 &
    reducedPartials_reducedPartials_36_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_385 = reducedPartials_reducedPartials_sum_384 ^ partials_36_15 ^
    partials_36_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_481 = reducedPartials_reducedPartials_sum_384 & partials_36_15 |
    partials_36_15 & partials_36_16 | reducedPartials_reducedPartials_sum_384 & partials_36_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_36_0_3 = reducedPartials_reducedPartials_sum_385 ^ partials_36_17 ^
    partials_36_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_482 = reducedPartials_reducedPartials_sum_385 & partials_36_17 |
    partials_36_17 & partials_36_18 | reducedPartials_reducedPartials_sum_385 & partials_36_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_386 = reducedPartials_reducedPartials_carry_482 ^
    reducedPartials_reducedPartials_carry_481 ^ reducedPartials_reducedPartials_carry_480; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_483 = reducedPartials_reducedPartials_carry_482 &
    reducedPartials_reducedPartials_carry_481 | reducedPartials_reducedPartials_carry_481 &
    reducedPartials_reducedPartials_carry_480 | reducedPartials_reducedPartials_carry_482 &
    reducedPartials_reducedPartials_carry_480; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_387 = reducedPartials_reducedPartials_sum_386 ^
    reducedPartials_reducedPartials_carry_479 ^ reducedPartials_reducedPartials_37_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_484 = reducedPartials_reducedPartials_sum_386 &
    reducedPartials_reducedPartials_carry_479 | reducedPartials_reducedPartials_carry_479 &
    reducedPartials_reducedPartials_37_0_1 | reducedPartials_reducedPartials_sum_386 &
    reducedPartials_reducedPartials_37_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_388 = reducedPartials_reducedPartials_sum_387 ^ partials_37_14 ^
    partials_37_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_485 = reducedPartials_reducedPartials_sum_387 & partials_37_14 |
    partials_37_14 & partials_37_15 | reducedPartials_reducedPartials_sum_387 & partials_37_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_37_0_2 = reducedPartials_reducedPartials_sum_388 ^ partials_37_16 ^
    partials_37_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_486 = reducedPartials_reducedPartials_sum_388 & partials_37_16 |
    partials_37_16 & partials_37_17 | reducedPartials_reducedPartials_sum_388 & partials_37_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_389 = reducedPartials_reducedPartials_carry_486 ^
    reducedPartials_reducedPartials_carry_485 ^ reducedPartials_reducedPartials_carry_484; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_487 = reducedPartials_reducedPartials_carry_486 &
    reducedPartials_reducedPartials_carry_485 | reducedPartials_reducedPartials_carry_485 &
    reducedPartials_reducedPartials_carry_484 | reducedPartials_reducedPartials_carry_486 &
    reducedPartials_reducedPartials_carry_484; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_390 = reducedPartials_reducedPartials_sum_389 ^
    reducedPartials_reducedPartials_carry_483 ^ reducedPartials_reducedPartials_38_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_488 = reducedPartials_reducedPartials_sum_389 &
    reducedPartials_reducedPartials_carry_483 | reducedPartials_reducedPartials_carry_483 &
    reducedPartials_reducedPartials_38_0_1 | reducedPartials_reducedPartials_sum_389 &
    reducedPartials_reducedPartials_38_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_391 = reducedPartials_reducedPartials_sum_390 ^ partials_38_13 ^
    partials_38_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_489 = reducedPartials_reducedPartials_sum_390 & partials_38_13 |
    partials_38_13 & partials_38_14 | reducedPartials_reducedPartials_sum_390 & partials_38_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_38_0_2 = reducedPartials_reducedPartials_sum_391 ^ partials_38_15 ^
    partials_38_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_490 = reducedPartials_reducedPartials_sum_391 & partials_38_15 |
    partials_38_15 & partials_38_16 | reducedPartials_reducedPartials_sum_391 & partials_38_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_392 = reducedPartials_reducedPartials_carry_490 ^
    reducedPartials_reducedPartials_carry_489 ^ reducedPartials_reducedPartials_carry_488; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_491 = reducedPartials_reducedPartials_carry_490 &
    reducedPartials_reducedPartials_carry_489 | reducedPartials_reducedPartials_carry_489 &
    reducedPartials_reducedPartials_carry_488 | reducedPartials_reducedPartials_carry_490 &
    reducedPartials_reducedPartials_carry_488; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_393 = reducedPartials_reducedPartials_sum_392 ^
    reducedPartials_reducedPartials_carry_487 ^ reducedPartials_reducedPartials_39_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_492 = reducedPartials_reducedPartials_sum_392 &
    reducedPartials_reducedPartials_carry_487 | reducedPartials_reducedPartials_carry_487 &
    reducedPartials_reducedPartials_39_0_1 | reducedPartials_reducedPartials_sum_392 &
    reducedPartials_reducedPartials_39_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_394 = reducedPartials_reducedPartials_sum_393 ^ partials_39_12 ^
    partials_39_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_493 = reducedPartials_reducedPartials_sum_393 & partials_39_12 |
    partials_39_12 & partials_39_13 | reducedPartials_reducedPartials_sum_393 & partials_39_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_39_0_2 = reducedPartials_reducedPartials_sum_394 ^ partials_39_14 ^
    partials_39_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_494 = reducedPartials_reducedPartials_sum_394 & partials_39_14 |
    partials_39_14 & partials_39_15 | reducedPartials_reducedPartials_sum_394 & partials_39_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_395 = reducedPartials_reducedPartials_carry_494 ^
    reducedPartials_reducedPartials_carry_493 ^ reducedPartials_reducedPartials_carry_492; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_495 = reducedPartials_reducedPartials_carry_494 &
    reducedPartials_reducedPartials_carry_493 | reducedPartials_reducedPartials_carry_493 &
    reducedPartials_reducedPartials_carry_492 | reducedPartials_reducedPartials_carry_494 &
    reducedPartials_reducedPartials_carry_492; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_396 = reducedPartials_reducedPartials_sum_395 ^
    reducedPartials_reducedPartials_carry_491 ^ reducedPartials_reducedPartials_40_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_496 = reducedPartials_reducedPartials_sum_395 &
    reducedPartials_reducedPartials_carry_491 | reducedPartials_reducedPartials_carry_491 &
    reducedPartials_reducedPartials_40_0_1 | reducedPartials_reducedPartials_sum_395 &
    reducedPartials_reducedPartials_40_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_397 = reducedPartials_reducedPartials_sum_396 ^ partials_40_11 ^
    partials_40_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_497 = reducedPartials_reducedPartials_sum_396 & partials_40_11 |
    partials_40_11 & partials_40_12 | reducedPartials_reducedPartials_sum_396 & partials_40_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_40_0_2 = reducedPartials_reducedPartials_sum_397 ^ partials_40_13 ^
    partials_40_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_498 = reducedPartials_reducedPartials_sum_397 & partials_40_13 |
    partials_40_13 & partials_40_14 | reducedPartials_reducedPartials_sum_397 & partials_40_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_398 = reducedPartials_reducedPartials_carry_498 ^
    reducedPartials_reducedPartials_carry_497 ^ reducedPartials_reducedPartials_carry_496; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_499 = reducedPartials_reducedPartials_carry_498 &
    reducedPartials_reducedPartials_carry_497 | reducedPartials_reducedPartials_carry_497 &
    reducedPartials_reducedPartials_carry_496 | reducedPartials_reducedPartials_carry_498 &
    reducedPartials_reducedPartials_carry_496; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_399 = reducedPartials_reducedPartials_sum_398 ^
    reducedPartials_reducedPartials_carry_495 ^ reducedPartials_reducedPartials_41_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_500 = reducedPartials_reducedPartials_sum_398 &
    reducedPartials_reducedPartials_carry_495 | reducedPartials_reducedPartials_carry_495 &
    reducedPartials_reducedPartials_41_0_1 | reducedPartials_reducedPartials_sum_398 &
    reducedPartials_reducedPartials_41_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_400 = reducedPartials_reducedPartials_sum_399 ^ partials_41_10 ^
    partials_41_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_501 = reducedPartials_reducedPartials_sum_399 & partials_41_10 |
    partials_41_10 & partials_41_11 | reducedPartials_reducedPartials_sum_399 & partials_41_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_41_0_2 = reducedPartials_reducedPartials_sum_400 ^ partials_41_12 ^
    partials_41_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_502 = reducedPartials_reducedPartials_sum_400 & partials_41_12 |
    partials_41_12 & partials_41_13 | reducedPartials_reducedPartials_sum_400 & partials_41_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_401 = reducedPartials_reducedPartials_carry_502 ^
    reducedPartials_reducedPartials_carry_501 ^ reducedPartials_reducedPartials_carry_500; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_503 = reducedPartials_reducedPartials_carry_502 &
    reducedPartials_reducedPartials_carry_501 | reducedPartials_reducedPartials_carry_501 &
    reducedPartials_reducedPartials_carry_500 | reducedPartials_reducedPartials_carry_502 &
    reducedPartials_reducedPartials_carry_500; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_402 = reducedPartials_reducedPartials_sum_401 ^
    reducedPartials_reducedPartials_carry_499 ^ reducedPartials_reducedPartials_42_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_504 = reducedPartials_reducedPartials_sum_401 &
    reducedPartials_reducedPartials_carry_499 | reducedPartials_reducedPartials_carry_499 &
    reducedPartials_reducedPartials_42_0_1 | reducedPartials_reducedPartials_sum_401 &
    reducedPartials_reducedPartials_42_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_403 = reducedPartials_reducedPartials_sum_402 ^ partials_42_9 ^
    partials_42_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_505 = reducedPartials_reducedPartials_sum_402 & partials_42_9 |
    partials_42_9 & partials_42_10 | reducedPartials_reducedPartials_sum_402 & partials_42_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_42_0_2 = reducedPartials_reducedPartials_sum_403 ^ partials_42_11 ^
    partials_42_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_506 = reducedPartials_reducedPartials_sum_403 & partials_42_11 |
    partials_42_11 & partials_42_12 | reducedPartials_reducedPartials_sum_403 & partials_42_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_404 = reducedPartials_reducedPartials_carry_506 ^
    reducedPartials_reducedPartials_carry_505 ^ reducedPartials_reducedPartials_carry_504; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_507 = reducedPartials_reducedPartials_carry_506 &
    reducedPartials_reducedPartials_carry_505 | reducedPartials_reducedPartials_carry_505 &
    reducedPartials_reducedPartials_carry_504 | reducedPartials_reducedPartials_carry_506 &
    reducedPartials_reducedPartials_carry_504; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_405 = reducedPartials_reducedPartials_sum_404 ^
    reducedPartials_reducedPartials_carry_503 ^ reducedPartials_reducedPartials_43_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_508 = reducedPartials_reducedPartials_sum_404 &
    reducedPartials_reducedPartials_carry_503 | reducedPartials_reducedPartials_carry_503 &
    reducedPartials_reducedPartials_43_0_1 | reducedPartials_reducedPartials_sum_404 &
    reducedPartials_reducedPartials_43_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_406 = reducedPartials_reducedPartials_sum_405 ^ partials_43_8 ^
    partials_43_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_509 = reducedPartials_reducedPartials_sum_405 & partials_43_8 |
    partials_43_8 & partials_43_9 | reducedPartials_reducedPartials_sum_405 & partials_43_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_43_0_2 = reducedPartials_reducedPartials_sum_406 ^ partials_43_10 ^
    partials_43_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_510 = reducedPartials_reducedPartials_sum_406 & partials_43_10 |
    partials_43_10 & partials_43_11 | reducedPartials_reducedPartials_sum_406 & partials_43_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_407 = reducedPartials_reducedPartials_carry_510 ^
    reducedPartials_reducedPartials_carry_509 ^ reducedPartials_reducedPartials_carry_508; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_511 = reducedPartials_reducedPartials_carry_510 &
    reducedPartials_reducedPartials_carry_509 | reducedPartials_reducedPartials_carry_509 &
    reducedPartials_reducedPartials_carry_508 | reducedPartials_reducedPartials_carry_510 &
    reducedPartials_reducedPartials_carry_508; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_408 = reducedPartials_reducedPartials_sum_407 ^
    reducedPartials_reducedPartials_carry_507 ^ reducedPartials_reducedPartials_44_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_512 = reducedPartials_reducedPartials_sum_407 &
    reducedPartials_reducedPartials_carry_507 | reducedPartials_reducedPartials_carry_507 &
    reducedPartials_reducedPartials_44_0_1 | reducedPartials_reducedPartials_sum_407 &
    reducedPartials_reducedPartials_44_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_409 = reducedPartials_reducedPartials_sum_408 ^ partials_44_7 ^
    partials_44_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_513 = reducedPartials_reducedPartials_sum_408 & partials_44_7 |
    partials_44_7 & partials_44_8 | reducedPartials_reducedPartials_sum_408 & partials_44_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_44_0_2 = reducedPartials_reducedPartials_sum_409 ^ partials_44_9 ^
    partials_44_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_514 = reducedPartials_reducedPartials_sum_409 & partials_44_9 |
    partials_44_9 & partials_44_10 | reducedPartials_reducedPartials_sum_409 & partials_44_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_410 = reducedPartials_reducedPartials_carry_514 ^
    reducedPartials_reducedPartials_carry_513 ^ reducedPartials_reducedPartials_carry_512; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_515 = reducedPartials_reducedPartials_carry_514 &
    reducedPartials_reducedPartials_carry_513 | reducedPartials_reducedPartials_carry_513 &
    reducedPartials_reducedPartials_carry_512 | reducedPartials_reducedPartials_carry_514 &
    reducedPartials_reducedPartials_carry_512; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_411 = reducedPartials_reducedPartials_sum_410 ^
    reducedPartials_reducedPartials_carry_511 ^ reducedPartials_reducedPartials_45_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_516 = reducedPartials_reducedPartials_sum_410 &
    reducedPartials_reducedPartials_carry_511 | reducedPartials_reducedPartials_carry_511 &
    reducedPartials_reducedPartials_45_0_1 | reducedPartials_reducedPartials_sum_410 &
    reducedPartials_reducedPartials_45_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_412 = reducedPartials_reducedPartials_sum_411 ^ partials_45_6 ^
    partials_45_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_517 = reducedPartials_reducedPartials_sum_411 & partials_45_6 |
    partials_45_6 & partials_45_7 | reducedPartials_reducedPartials_sum_411 & partials_45_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_45_0_2 = reducedPartials_reducedPartials_sum_412 ^ partials_45_8 ^ partials_45_9
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_518 = reducedPartials_reducedPartials_sum_412 & partials_45_8 |
    partials_45_8 & partials_45_9 | reducedPartials_reducedPartials_sum_412 & partials_45_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_413 = reducedPartials_reducedPartials_carry_518 ^
    reducedPartials_reducedPartials_carry_517 ^ reducedPartials_reducedPartials_carry_516; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_519 = reducedPartials_reducedPartials_carry_518 &
    reducedPartials_reducedPartials_carry_517 | reducedPartials_reducedPartials_carry_517 &
    reducedPartials_reducedPartials_carry_516 | reducedPartials_reducedPartials_carry_518 &
    reducedPartials_reducedPartials_carry_516; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_414 = reducedPartials_reducedPartials_sum_413 ^
    reducedPartials_reducedPartials_carry_515 ^ reducedPartials_reducedPartials_46_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_520 = reducedPartials_reducedPartials_sum_413 &
    reducedPartials_reducedPartials_carry_515 | reducedPartials_reducedPartials_carry_515 &
    reducedPartials_reducedPartials_46_0 | reducedPartials_reducedPartials_sum_413 &
    reducedPartials_reducedPartials_46_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_415 = reducedPartials_reducedPartials_sum_414 ^ partials_46_5 ^
    partials_46_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_521 = reducedPartials_reducedPartials_sum_414 & partials_46_5 |
    partials_46_5 & partials_46_6 | reducedPartials_reducedPartials_sum_414 & partials_46_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_46_0_1 = reducedPartials_reducedPartials_sum_415 ^ partials_46_7 ^ partials_46_8
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_522 = reducedPartials_reducedPartials_sum_415 & partials_46_7 |
    partials_46_7 & partials_46_8 | reducedPartials_reducedPartials_sum_415 & partials_46_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_416 = reducedPartials_reducedPartials_carry_522 ^
    reducedPartials_reducedPartials_carry_521 ^ reducedPartials_reducedPartials_carry_520; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_523 = reducedPartials_reducedPartials_carry_522 &
    reducedPartials_reducedPartials_carry_521 | reducedPartials_reducedPartials_carry_521 &
    reducedPartials_reducedPartials_carry_520 | reducedPartials_reducedPartials_carry_522 &
    reducedPartials_reducedPartials_carry_520; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_417 = reducedPartials_reducedPartials_sum_416 ^
    reducedPartials_reducedPartials_carry_519 ^ reducedPartials_reducedPartials_47_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_524 = reducedPartials_reducedPartials_sum_416 &
    reducedPartials_reducedPartials_carry_519 | reducedPartials_reducedPartials_carry_519 &
    reducedPartials_reducedPartials_47_0 | reducedPartials_reducedPartials_sum_416 &
    reducedPartials_reducedPartials_47_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_418 = reducedPartials_reducedPartials_sum_417 ^ partials_47_4 ^
    partials_47_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_525 = reducedPartials_reducedPartials_sum_417 & partials_47_4 |
    partials_47_4 & partials_47_5 | reducedPartials_reducedPartials_sum_417 & partials_47_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_47_0_1 = reducedPartials_reducedPartials_sum_418 ^ partials_47_6 ^ partials_47_7
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_526 = reducedPartials_reducedPartials_sum_418 & partials_47_6 |
    partials_47_6 & partials_47_7 | reducedPartials_reducedPartials_sum_418 & partials_47_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_419 = reducedPartials_reducedPartials_carry_526 ^
    reducedPartials_reducedPartials_carry_525 ^ reducedPartials_reducedPartials_carry_524; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_527 = reducedPartials_reducedPartials_carry_526 &
    reducedPartials_reducedPartials_carry_525 | reducedPartials_reducedPartials_carry_525 &
    reducedPartials_reducedPartials_carry_524 | reducedPartials_reducedPartials_carry_526 &
    reducedPartials_reducedPartials_carry_524; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_420 = reducedPartials_reducedPartials_sum_419 ^
    reducedPartials_reducedPartials_carry_523 ^ reducedPartials_reducedPartials_48_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_528 = reducedPartials_reducedPartials_sum_419 &
    reducedPartials_reducedPartials_carry_523 | reducedPartials_reducedPartials_carry_523 &
    reducedPartials_reducedPartials_48_0 | reducedPartials_reducedPartials_sum_419 &
    reducedPartials_reducedPartials_48_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_421 = reducedPartials_reducedPartials_sum_420 ^ partials_48_3 ^
    partials_48_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_529 = reducedPartials_reducedPartials_sum_420 & partials_48_3 |
    partials_48_3 & partials_48_4 | reducedPartials_reducedPartials_sum_420 & partials_48_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_48_0_1 = reducedPartials_reducedPartials_sum_421 ^ partials_48_5 ^ partials_48_6
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_530 = reducedPartials_reducedPartials_sum_421 & partials_48_5 |
    partials_48_5 & partials_48_6 | reducedPartials_reducedPartials_sum_421 & partials_48_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_422 = reducedPartials_reducedPartials_carry_530 ^
    reducedPartials_reducedPartials_carry_529 ^ reducedPartials_reducedPartials_carry_528; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_531 = reducedPartials_reducedPartials_carry_530 &
    reducedPartials_reducedPartials_carry_529 | reducedPartials_reducedPartials_carry_529 &
    reducedPartials_reducedPartials_carry_528 | reducedPartials_reducedPartials_carry_530 &
    reducedPartials_reducedPartials_carry_528; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_423 = reducedPartials_reducedPartials_sum_422 ^
    reducedPartials_reducedPartials_carry_527 ^ reducedPartials_reducedPartials_49_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_532 = reducedPartials_reducedPartials_sum_422 &
    reducedPartials_reducedPartials_carry_527 | reducedPartials_reducedPartials_carry_527 &
    reducedPartials_reducedPartials_49_0 | reducedPartials_reducedPartials_sum_422 &
    reducedPartials_reducedPartials_49_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_424 = reducedPartials_reducedPartials_sum_423 ^ partials_49_2 ^
    partials_49_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_533 = reducedPartials_reducedPartials_sum_423 & partials_49_2 |
    partials_49_2 & partials_49_3 | reducedPartials_reducedPartials_sum_423 & partials_49_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_49_0_1 = reducedPartials_reducedPartials_sum_424 ^ partials_49_4 ^ partials_49_5
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_534 = reducedPartials_reducedPartials_sum_424 & partials_49_4 |
    partials_49_4 & partials_49_5 | reducedPartials_reducedPartials_sum_424 & partials_49_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_425 = reducedPartials_reducedPartials_carry_534 ^
    reducedPartials_reducedPartials_carry_533 ^ reducedPartials_reducedPartials_carry_532; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_535 = reducedPartials_reducedPartials_carry_534 &
    reducedPartials_reducedPartials_carry_533 | reducedPartials_reducedPartials_carry_533 &
    reducedPartials_reducedPartials_carry_532 | reducedPartials_reducedPartials_carry_534 &
    reducedPartials_reducedPartials_carry_532; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_426 = reducedPartials_reducedPartials_sum_425 ^
    reducedPartials_reducedPartials_carry_531 ^ reducedPartials_reducedPartials_50_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_536 = reducedPartials_reducedPartials_sum_425 &
    reducedPartials_reducedPartials_carry_531 | reducedPartials_reducedPartials_carry_531 &
    reducedPartials_reducedPartials_50_0 | reducedPartials_reducedPartials_sum_425 &
    reducedPartials_reducedPartials_50_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_427 = reducedPartials_reducedPartials_sum_426 ^ partials_50_1 ^
    partials_50_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_537 = reducedPartials_reducedPartials_sum_426 & partials_50_1 |
    partials_50_1 & partials_50_2 | reducedPartials_reducedPartials_sum_426 & partials_50_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_50_0_1 = reducedPartials_reducedPartials_sum_427 ^ partials_50_3 ^ partials_50_4
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_538 = reducedPartials_reducedPartials_sum_427 & partials_50_3 |
    partials_50_3 & partials_50_4 | reducedPartials_reducedPartials_sum_427 & partials_50_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_428 = reducedPartials_reducedPartials_carry_538 ^
    reducedPartials_reducedPartials_carry_537 ^ reducedPartials_reducedPartials_carry_536; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_539 = reducedPartials_reducedPartials_carry_538 &
    reducedPartials_reducedPartials_carry_537 | reducedPartials_reducedPartials_carry_537 &
    reducedPartials_reducedPartials_carry_536 | reducedPartials_reducedPartials_carry_538 &
    reducedPartials_reducedPartials_carry_536; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_429 = reducedPartials_reducedPartials_sum_428 ^
    reducedPartials_reducedPartials_carry_535 ^ reducedPartials_reducedPartials_51_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_540 = reducedPartials_reducedPartials_sum_428 &
    reducedPartials_reducedPartials_carry_535 | reducedPartials_reducedPartials_carry_535 &
    reducedPartials_reducedPartials_51_0 | reducedPartials_reducedPartials_sum_428 &
    reducedPartials_reducedPartials_51_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_430 = reducedPartials_reducedPartials_sum_429 ^ partials_51_0 ^
    partials_51_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_541 = reducedPartials_reducedPartials_sum_429 & partials_51_0 |
    partials_51_0 & partials_51_1 | reducedPartials_reducedPartials_sum_429 & partials_51_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_51_0_1 = reducedPartials_reducedPartials_sum_430 ^ partials_51_2 ^ partials_51_3
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_542 = reducedPartials_reducedPartials_sum_430 & partials_51_2 |
    partials_51_2 & partials_51_3 | reducedPartials_reducedPartials_sum_430 & partials_51_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_431 = reducedPartials_reducedPartials_carry_542 ^
    reducedPartials_reducedPartials_carry_541 ^ reducedPartials_reducedPartials_carry_540; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_543 = reducedPartials_reducedPartials_carry_542 &
    reducedPartials_reducedPartials_carry_541 | reducedPartials_reducedPartials_carry_541 &
    reducedPartials_reducedPartials_carry_540 | reducedPartials_reducedPartials_carry_542 &
    reducedPartials_reducedPartials_carry_540; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_432 = reducedPartials_reducedPartials_sum_431 ^
    reducedPartials_reducedPartials_carry_539 ^ partials_52_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_544 = reducedPartials_reducedPartials_sum_431 &
    reducedPartials_reducedPartials_carry_539 | reducedPartials_reducedPartials_carry_539 & partials_52_0 |
    reducedPartials_reducedPartials_sum_431 & partials_52_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_52_0 = reducedPartials_reducedPartials_sum_432 ^ partials_52_1 ^ partials_52_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_545 = reducedPartials_reducedPartials_sum_432 & partials_52_1 |
    partials_52_1 & partials_52_2 | reducedPartials_reducedPartials_sum_432 & partials_52_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_433 = reducedPartials_reducedPartials_carry_545 ^
    reducedPartials_reducedPartials_carry_544 ^ reducedPartials_reducedPartials_carry_543; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_546 = reducedPartials_reducedPartials_carry_545 &
    reducedPartials_reducedPartials_carry_544 | reducedPartials_reducedPartials_carry_544 &
    reducedPartials_reducedPartials_carry_543 | reducedPartials_reducedPartials_carry_545 &
    reducedPartials_reducedPartials_carry_543; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_53_0 = reducedPartials_reducedPartials_sum_433 ^ partials_53_0 ^ partials_53_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_547 = reducedPartials_reducedPartials_sum_433 & partials_53_0 |
    partials_53_0 & partials_53_1 | reducedPartials_reducedPartials_sum_433 & partials_53_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_54_0 = reducedPartials_reducedPartials_carry_547 ^
    reducedPartials_reducedPartials_carry_546 ^ partials_54_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_55_0 = reducedPartials_reducedPartials_carry_547 &
    reducedPartials_reducedPartials_carry_546 | reducedPartials_reducedPartials_carry_546 & partials_54_0 |
    reducedPartials_reducedPartials_carry_547 & partials_54_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_6_0 = partials_6_0 ^ partials_6_1; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_548 = partials_6_0 & partials_6_1; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_434 = reducedPartials_reducedPartials_carry_548 ^ partials_7_0 ^
    partials_7_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_549 = reducedPartials_reducedPartials_carry_548 & partials_7_0 |
    partials_7_0 & partials_7_1 | reducedPartials_reducedPartials_carry_548 & partials_7_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_7_0 = reducedPartials_reducedPartials_sum_434 ^ partials_7_2; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_550 = reducedPartials_reducedPartials_sum_434 & partials_7_2; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_435 = reducedPartials_reducedPartials_carry_550 ^
    reducedPartials_reducedPartials_carry_549 ^ partials_8_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_551 = reducedPartials_reducedPartials_carry_550 &
    reducedPartials_reducedPartials_carry_549 | reducedPartials_reducedPartials_carry_549 & partials_8_0 |
    reducedPartials_reducedPartials_carry_550 & partials_8_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_436 = reducedPartials_reducedPartials_sum_435 ^ partials_8_1 ^ partials_8_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_552 = reducedPartials_reducedPartials_sum_435 & partials_8_1 |
    partials_8_1 & partials_8_2 | reducedPartials_reducedPartials_sum_435 & partials_8_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_8_0 = reducedPartials_reducedPartials_sum_436 ^ partials_8_3; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_553 = reducedPartials_reducedPartials_sum_436 & partials_8_3; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_437 = reducedPartials_reducedPartials_carry_553 ^
    reducedPartials_reducedPartials_carry_552 ^ reducedPartials_reducedPartials_carry_551; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_554 = reducedPartials_reducedPartials_carry_553 &
    reducedPartials_reducedPartials_carry_552 | reducedPartials_reducedPartials_carry_552 &
    reducedPartials_reducedPartials_carry_551 | reducedPartials_reducedPartials_carry_553 &
    reducedPartials_reducedPartials_carry_551; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_438 = reducedPartials_reducedPartials_sum_437 ^
    reducedPartials_reducedPartials_9_0 ^ partials_9_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_555 = reducedPartials_reducedPartials_sum_437 &
    reducedPartials_reducedPartials_9_0 | reducedPartials_reducedPartials_9_0 & partials_9_2 |
    reducedPartials_reducedPartials_sum_437 & partials_9_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_9_0_1 = reducedPartials_reducedPartials_sum_438 ^ partials_9_3 ^ partials_9_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_556 = reducedPartials_reducedPartials_sum_438 & partials_9_3 |
    partials_9_3 & partials_9_4 | reducedPartials_reducedPartials_sum_438 & partials_9_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_439 = reducedPartials_reducedPartials_carry_556 ^
    reducedPartials_reducedPartials_carry_555 ^ reducedPartials_reducedPartials_carry_554; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_557 = reducedPartials_reducedPartials_carry_556 &
    reducedPartials_reducedPartials_carry_555 | reducedPartials_reducedPartials_carry_555 &
    reducedPartials_reducedPartials_carry_554 | reducedPartials_reducedPartials_carry_556 &
    reducedPartials_reducedPartials_carry_554; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_440 = reducedPartials_reducedPartials_sum_439 ^
    reducedPartials_reducedPartials_10_0 ^ partials_10_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_558 = reducedPartials_reducedPartials_sum_439 &
    reducedPartials_reducedPartials_10_0 | reducedPartials_reducedPartials_10_0 & partials_10_3 |
    reducedPartials_reducedPartials_sum_439 & partials_10_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_10_0_1 = reducedPartials_reducedPartials_sum_440 ^ partials_10_4 ^ partials_10_5
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_559 = reducedPartials_reducedPartials_sum_440 & partials_10_4 |
    partials_10_4 & partials_10_5 | reducedPartials_reducedPartials_sum_440 & partials_10_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_441 = reducedPartials_reducedPartials_carry_559 ^
    reducedPartials_reducedPartials_carry_558 ^ reducedPartials_reducedPartials_carry_557; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_560 = reducedPartials_reducedPartials_carry_559 &
    reducedPartials_reducedPartials_carry_558 | reducedPartials_reducedPartials_carry_558 &
    reducedPartials_reducedPartials_carry_557 | reducedPartials_reducedPartials_carry_559 &
    reducedPartials_reducedPartials_carry_557; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_442 = reducedPartials_reducedPartials_sum_441 ^
    reducedPartials_reducedPartials_11_0 ^ partials_11_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_561 = reducedPartials_reducedPartials_sum_441 &
    reducedPartials_reducedPartials_11_0 | reducedPartials_reducedPartials_11_0 & partials_11_4 |
    reducedPartials_reducedPartials_sum_441 & partials_11_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_11_0_1 = reducedPartials_reducedPartials_sum_442 ^ partials_11_5 ^ partials_11_6
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_562 = reducedPartials_reducedPartials_sum_442 & partials_11_5 |
    partials_11_5 & partials_11_6 | reducedPartials_reducedPartials_sum_442 & partials_11_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_443 = reducedPartials_reducedPartials_carry_562 ^
    reducedPartials_reducedPartials_carry_561 ^ reducedPartials_reducedPartials_carry_560; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_563 = reducedPartials_reducedPartials_carry_562 &
    reducedPartials_reducedPartials_carry_561 | reducedPartials_reducedPartials_carry_561 &
    reducedPartials_reducedPartials_carry_560 | reducedPartials_reducedPartials_carry_562 &
    reducedPartials_reducedPartials_carry_560; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_444 = reducedPartials_reducedPartials_sum_443 ^
    reducedPartials_reducedPartials_12_0 ^ partials_12_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_564 = reducedPartials_reducedPartials_sum_443 &
    reducedPartials_reducedPartials_12_0 | reducedPartials_reducedPartials_12_0 & partials_12_5 |
    reducedPartials_reducedPartials_sum_443 & partials_12_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_12_0_1 = reducedPartials_reducedPartials_sum_444 ^ partials_12_6 ^ partials_12_7
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_565 = reducedPartials_reducedPartials_sum_444 & partials_12_6 |
    partials_12_6 & partials_12_7 | reducedPartials_reducedPartials_sum_444 & partials_12_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_445 = reducedPartials_reducedPartials_carry_565 ^
    reducedPartials_reducedPartials_carry_564 ^ reducedPartials_reducedPartials_carry_563; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_566 = reducedPartials_reducedPartials_carry_565 &
    reducedPartials_reducedPartials_carry_564 | reducedPartials_reducedPartials_carry_564 &
    reducedPartials_reducedPartials_carry_563 | reducedPartials_reducedPartials_carry_565 &
    reducedPartials_reducedPartials_carry_563; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_446 = reducedPartials_reducedPartials_sum_445 ^
    reducedPartials_reducedPartials_13_0_1 ^ partials_13_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_567 = reducedPartials_reducedPartials_sum_445 &
    reducedPartials_reducedPartials_13_0_1 | reducedPartials_reducedPartials_13_0_1 & partials_13_6 |
    reducedPartials_reducedPartials_sum_445 & partials_13_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_13_0_2 = reducedPartials_reducedPartials_sum_446 ^ partials_13_7 ^ partials_13_8
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_568 = reducedPartials_reducedPartials_sum_446 & partials_13_7 |
    partials_13_7 & partials_13_8 | reducedPartials_reducedPartials_sum_446 & partials_13_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_447 = reducedPartials_reducedPartials_carry_568 ^
    reducedPartials_reducedPartials_carry_567 ^ reducedPartials_reducedPartials_carry_566; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_569 = reducedPartials_reducedPartials_carry_568 &
    reducedPartials_reducedPartials_carry_567 | reducedPartials_reducedPartials_carry_567 &
    reducedPartials_reducedPartials_carry_566 | reducedPartials_reducedPartials_carry_568 &
    reducedPartials_reducedPartials_carry_566; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_448 = reducedPartials_reducedPartials_sum_447 ^
    reducedPartials_reducedPartials_14_0_1 ^ partials_14_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_570 = reducedPartials_reducedPartials_sum_447 &
    reducedPartials_reducedPartials_14_0_1 | reducedPartials_reducedPartials_14_0_1 & partials_14_7 |
    reducedPartials_reducedPartials_sum_447 & partials_14_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_14_0_2 = reducedPartials_reducedPartials_sum_448 ^ partials_14_8 ^ partials_14_9
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_571 = reducedPartials_reducedPartials_sum_448 & partials_14_8 |
    partials_14_8 & partials_14_9 | reducedPartials_reducedPartials_sum_448 & partials_14_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_449 = reducedPartials_reducedPartials_carry_571 ^
    reducedPartials_reducedPartials_carry_570 ^ reducedPartials_reducedPartials_carry_569; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_572 = reducedPartials_reducedPartials_carry_571 &
    reducedPartials_reducedPartials_carry_570 | reducedPartials_reducedPartials_carry_570 &
    reducedPartials_reducedPartials_carry_569 | reducedPartials_reducedPartials_carry_571 &
    reducedPartials_reducedPartials_carry_569; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_450 = reducedPartials_reducedPartials_sum_449 ^
    reducedPartials_reducedPartials_15_0_1 ^ partials_15_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_573 = reducedPartials_reducedPartials_sum_449 &
    reducedPartials_reducedPartials_15_0_1 | reducedPartials_reducedPartials_15_0_1 & partials_15_8 |
    reducedPartials_reducedPartials_sum_449 & partials_15_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_15_0_2 = reducedPartials_reducedPartials_sum_450 ^ partials_15_9 ^
    partials_15_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_574 = reducedPartials_reducedPartials_sum_450 & partials_15_9 |
    partials_15_9 & partials_15_10 | reducedPartials_reducedPartials_sum_450 & partials_15_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_451 = reducedPartials_reducedPartials_carry_574 ^
    reducedPartials_reducedPartials_carry_573 ^ reducedPartials_reducedPartials_carry_572; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_575 = reducedPartials_reducedPartials_carry_574 &
    reducedPartials_reducedPartials_carry_573 | reducedPartials_reducedPartials_carry_573 &
    reducedPartials_reducedPartials_carry_572 | reducedPartials_reducedPartials_carry_574 &
    reducedPartials_reducedPartials_carry_572; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_452 = reducedPartials_reducedPartials_sum_451 ^
    reducedPartials_reducedPartials_16_0_1 ^ partials_16_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_576 = reducedPartials_reducedPartials_sum_451 &
    reducedPartials_reducedPartials_16_0_1 | reducedPartials_reducedPartials_16_0_1 & partials_16_9 |
    reducedPartials_reducedPartials_sum_451 & partials_16_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_16_0_2 = reducedPartials_reducedPartials_sum_452 ^ partials_16_10 ^
    partials_16_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_577 = reducedPartials_reducedPartials_sum_452 & partials_16_10 |
    partials_16_10 & partials_16_11 | reducedPartials_reducedPartials_sum_452 & partials_16_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_453 = reducedPartials_reducedPartials_carry_577 ^
    reducedPartials_reducedPartials_carry_576 ^ reducedPartials_reducedPartials_carry_575; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_578 = reducedPartials_reducedPartials_carry_577 &
    reducedPartials_reducedPartials_carry_576 | reducedPartials_reducedPartials_carry_576 &
    reducedPartials_reducedPartials_carry_575 | reducedPartials_reducedPartials_carry_577 &
    reducedPartials_reducedPartials_carry_575; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_454 = reducedPartials_reducedPartials_sum_453 ^
    reducedPartials_reducedPartials_17_0_1 ^ partials_17_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_579 = reducedPartials_reducedPartials_sum_453 &
    reducedPartials_reducedPartials_17_0_1 | reducedPartials_reducedPartials_17_0_1 & partials_17_10 |
    reducedPartials_reducedPartials_sum_453 & partials_17_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_17_0_2 = reducedPartials_reducedPartials_sum_454 ^ partials_17_11 ^
    partials_17_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_580 = reducedPartials_reducedPartials_sum_454 & partials_17_11 |
    partials_17_11 & partials_17_12 | reducedPartials_reducedPartials_sum_454 & partials_17_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_455 = reducedPartials_reducedPartials_carry_580 ^
    reducedPartials_reducedPartials_carry_579 ^ reducedPartials_reducedPartials_carry_578; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_581 = reducedPartials_reducedPartials_carry_580 &
    reducedPartials_reducedPartials_carry_579 | reducedPartials_reducedPartials_carry_579 &
    reducedPartials_reducedPartials_carry_578 | reducedPartials_reducedPartials_carry_580 &
    reducedPartials_reducedPartials_carry_578; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_456 = reducedPartials_reducedPartials_sum_455 ^
    reducedPartials_reducedPartials_18_0_1 ^ partials_18_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_582 = reducedPartials_reducedPartials_sum_455 &
    reducedPartials_reducedPartials_18_0_1 | reducedPartials_reducedPartials_18_0_1 & partials_18_11 |
    reducedPartials_reducedPartials_sum_455 & partials_18_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_18_0_2 = reducedPartials_reducedPartials_sum_456 ^ partials_18_12 ^
    partials_18_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_583 = reducedPartials_reducedPartials_sum_456 & partials_18_12 |
    partials_18_12 & partials_18_13 | reducedPartials_reducedPartials_sum_456 & partials_18_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_457 = reducedPartials_reducedPartials_carry_583 ^
    reducedPartials_reducedPartials_carry_582 ^ reducedPartials_reducedPartials_carry_581; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_584 = reducedPartials_reducedPartials_carry_583 &
    reducedPartials_reducedPartials_carry_582 | reducedPartials_reducedPartials_carry_582 &
    reducedPartials_reducedPartials_carry_581 | reducedPartials_reducedPartials_carry_583 &
    reducedPartials_reducedPartials_carry_581; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_458 = reducedPartials_reducedPartials_sum_457 ^
    reducedPartials_reducedPartials_19_0_2 ^ partials_19_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_585 = reducedPartials_reducedPartials_sum_457 &
    reducedPartials_reducedPartials_19_0_2 | reducedPartials_reducedPartials_19_0_2 & partials_19_12 |
    reducedPartials_reducedPartials_sum_457 & partials_19_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_19_0_3 = reducedPartials_reducedPartials_sum_458 ^ partials_19_13 ^
    partials_19_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_586 = reducedPartials_reducedPartials_sum_458 & partials_19_13 |
    partials_19_13 & partials_19_14 | reducedPartials_reducedPartials_sum_458 & partials_19_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_459 = reducedPartials_reducedPartials_carry_586 ^
    reducedPartials_reducedPartials_carry_585 ^ reducedPartials_reducedPartials_carry_584; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_587 = reducedPartials_reducedPartials_carry_586 &
    reducedPartials_reducedPartials_carry_585 | reducedPartials_reducedPartials_carry_585 &
    reducedPartials_reducedPartials_carry_584 | reducedPartials_reducedPartials_carry_586 &
    reducedPartials_reducedPartials_carry_584; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_460 = reducedPartials_reducedPartials_sum_459 ^
    reducedPartials_reducedPartials_20_0_2 ^ partials_20_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_588 = reducedPartials_reducedPartials_sum_459 &
    reducedPartials_reducedPartials_20_0_2 | reducedPartials_reducedPartials_20_0_2 & partials_20_13 |
    reducedPartials_reducedPartials_sum_459 & partials_20_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_20_0_3 = reducedPartials_reducedPartials_sum_460 ^ partials_20_14 ^
    partials_20_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_589 = reducedPartials_reducedPartials_sum_460 & partials_20_14 |
    partials_20_14 & partials_20_15 | reducedPartials_reducedPartials_sum_460 & partials_20_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_461 = reducedPartials_reducedPartials_carry_589 ^
    reducedPartials_reducedPartials_carry_588 ^ reducedPartials_reducedPartials_carry_587; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_590 = reducedPartials_reducedPartials_carry_589 &
    reducedPartials_reducedPartials_carry_588 | reducedPartials_reducedPartials_carry_588 &
    reducedPartials_reducedPartials_carry_587 | reducedPartials_reducedPartials_carry_589 &
    reducedPartials_reducedPartials_carry_587; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_462 = reducedPartials_reducedPartials_sum_461 ^
    reducedPartials_reducedPartials_21_0_2 ^ partials_21_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_591 = reducedPartials_reducedPartials_sum_461 &
    reducedPartials_reducedPartials_21_0_2 | reducedPartials_reducedPartials_21_0_2 & partials_21_14 |
    reducedPartials_reducedPartials_sum_461 & partials_21_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_21_0_3 = reducedPartials_reducedPartials_sum_462 ^ partials_21_15 ^
    partials_21_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_592 = reducedPartials_reducedPartials_sum_462 & partials_21_15 |
    partials_21_15 & partials_21_16 | reducedPartials_reducedPartials_sum_462 & partials_21_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_463 = reducedPartials_reducedPartials_carry_592 ^
    reducedPartials_reducedPartials_carry_591 ^ reducedPartials_reducedPartials_carry_590; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_593 = reducedPartials_reducedPartials_carry_592 &
    reducedPartials_reducedPartials_carry_591 | reducedPartials_reducedPartials_carry_591 &
    reducedPartials_reducedPartials_carry_590 | reducedPartials_reducedPartials_carry_592 &
    reducedPartials_reducedPartials_carry_590; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_464 = reducedPartials_reducedPartials_sum_463 ^
    reducedPartials_reducedPartials_22_0_2 ^ partials_22_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_594 = reducedPartials_reducedPartials_sum_463 &
    reducedPartials_reducedPartials_22_0_2 | reducedPartials_reducedPartials_22_0_2 & partials_22_15 |
    reducedPartials_reducedPartials_sum_463 & partials_22_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_22_0_3 = reducedPartials_reducedPartials_sum_464 ^ partials_22_16 ^
    partials_22_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_595 = reducedPartials_reducedPartials_sum_464 & partials_22_16 |
    partials_22_16 & partials_22_17 | reducedPartials_reducedPartials_sum_464 & partials_22_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_465 = reducedPartials_reducedPartials_carry_595 ^
    reducedPartials_reducedPartials_carry_594 ^ reducedPartials_reducedPartials_carry_593; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_596 = reducedPartials_reducedPartials_carry_595 &
    reducedPartials_reducedPartials_carry_594 | reducedPartials_reducedPartials_carry_594 &
    reducedPartials_reducedPartials_carry_593 | reducedPartials_reducedPartials_carry_595 &
    reducedPartials_reducedPartials_carry_593; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_466 = reducedPartials_reducedPartials_sum_465 ^
    reducedPartials_reducedPartials_23_0_2 ^ partials_23_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_597 = reducedPartials_reducedPartials_sum_465 &
    reducedPartials_reducedPartials_23_0_2 | reducedPartials_reducedPartials_23_0_2 & partials_23_16 |
    reducedPartials_reducedPartials_sum_465 & partials_23_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_23_0_3 = reducedPartials_reducedPartials_sum_466 ^ partials_23_17 ^
    partials_23_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_598 = reducedPartials_reducedPartials_sum_466 & partials_23_17 |
    partials_23_17 & partials_23_18 | reducedPartials_reducedPartials_sum_466 & partials_23_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_467 = reducedPartials_reducedPartials_carry_598 ^
    reducedPartials_reducedPartials_carry_597 ^ reducedPartials_reducedPartials_carry_596; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_599 = reducedPartials_reducedPartials_carry_598 &
    reducedPartials_reducedPartials_carry_597 | reducedPartials_reducedPartials_carry_597 &
    reducedPartials_reducedPartials_carry_596 | reducedPartials_reducedPartials_carry_598 &
    reducedPartials_reducedPartials_carry_596; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_468 = reducedPartials_reducedPartials_sum_467 ^
    reducedPartials_reducedPartials_24_0_2 ^ partials_24_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_600 = reducedPartials_reducedPartials_sum_467 &
    reducedPartials_reducedPartials_24_0_2 | reducedPartials_reducedPartials_24_0_2 & partials_24_17 |
    reducedPartials_reducedPartials_sum_467 & partials_24_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_24_0_3 = reducedPartials_reducedPartials_sum_468 ^ partials_24_18 ^
    partials_24_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_601 = reducedPartials_reducedPartials_sum_468 & partials_24_18 |
    partials_24_18 & partials_24_19 | reducedPartials_reducedPartials_sum_468 & partials_24_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_469 = reducedPartials_reducedPartials_carry_601 ^
    reducedPartials_reducedPartials_carry_600 ^ reducedPartials_reducedPartials_carry_599; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_602 = reducedPartials_reducedPartials_carry_601 &
    reducedPartials_reducedPartials_carry_600 | reducedPartials_reducedPartials_carry_600 &
    reducedPartials_reducedPartials_carry_599 | reducedPartials_reducedPartials_carry_601 &
    reducedPartials_reducedPartials_carry_599; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_470 = reducedPartials_reducedPartials_sum_469 ^
    reducedPartials_reducedPartials_25_0_2 ^ partials_25_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_603 = reducedPartials_reducedPartials_sum_469 &
    reducedPartials_reducedPartials_25_0_2 | reducedPartials_reducedPartials_25_0_2 & partials_25_18 |
    reducedPartials_reducedPartials_sum_469 & partials_25_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_25_0_3 = reducedPartials_reducedPartials_sum_470 ^ partials_25_19 ^
    partials_25_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_604 = reducedPartials_reducedPartials_sum_470 & partials_25_19 |
    partials_25_19 & partials_25_20 | reducedPartials_reducedPartials_sum_470 & partials_25_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_471 = reducedPartials_reducedPartials_carry_604 ^
    reducedPartials_reducedPartials_carry_603 ^ reducedPartials_reducedPartials_carry_602; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_605 = reducedPartials_reducedPartials_carry_604 &
    reducedPartials_reducedPartials_carry_603 | reducedPartials_reducedPartials_carry_603 &
    reducedPartials_reducedPartials_carry_602 | reducedPartials_reducedPartials_carry_604 &
    reducedPartials_reducedPartials_carry_602; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_472 = reducedPartials_reducedPartials_sum_471 ^
    reducedPartials_reducedPartials_26_0_2 ^ partials_26_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_606 = reducedPartials_reducedPartials_sum_471 &
    reducedPartials_reducedPartials_26_0_2 | reducedPartials_reducedPartials_26_0_2 & partials_26_19 |
    reducedPartials_reducedPartials_sum_471 & partials_26_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_26_0_3 = reducedPartials_reducedPartials_sum_472 ^ partials_26_20 ^
    partials_26_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_607 = reducedPartials_reducedPartials_sum_472 & partials_26_20 |
    partials_26_20 & partials_26_21 | reducedPartials_reducedPartials_sum_472 & partials_26_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_473 = reducedPartials_reducedPartials_carry_607 ^
    reducedPartials_reducedPartials_carry_606 ^ reducedPartials_reducedPartials_carry_605; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_608 = reducedPartials_reducedPartials_carry_607 &
    reducedPartials_reducedPartials_carry_606 | reducedPartials_reducedPartials_carry_606 &
    reducedPartials_reducedPartials_carry_605 | reducedPartials_reducedPartials_carry_607 &
    reducedPartials_reducedPartials_carry_605; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_474 = reducedPartials_reducedPartials_sum_473 ^
    reducedPartials_reducedPartials_27_0_2 ^ partials_27_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_609 = reducedPartials_reducedPartials_sum_473 &
    reducedPartials_reducedPartials_27_0_2 | reducedPartials_reducedPartials_27_0_2 & partials_27_20 |
    reducedPartials_reducedPartials_sum_473 & partials_27_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_27_0_3 = reducedPartials_reducedPartials_sum_474 ^ partials_27_21 ^
    partials_27_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_610 = reducedPartials_reducedPartials_sum_474 & partials_27_21 |
    partials_27_21 & partials_27_22 | reducedPartials_reducedPartials_sum_474 & partials_27_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_475 = reducedPartials_reducedPartials_carry_610 ^
    reducedPartials_reducedPartials_carry_609 ^ reducedPartials_reducedPartials_carry_608; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_611 = reducedPartials_reducedPartials_carry_610 &
    reducedPartials_reducedPartials_carry_609 | reducedPartials_reducedPartials_carry_609 &
    reducedPartials_reducedPartials_carry_608 | reducedPartials_reducedPartials_carry_610 &
    reducedPartials_reducedPartials_carry_608; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_476 = reducedPartials_reducedPartials_sum_475 ^
    reducedPartials_reducedPartials_28_0_3 ^ partials_28_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_612 = reducedPartials_reducedPartials_sum_475 &
    reducedPartials_reducedPartials_28_0_3 | reducedPartials_reducedPartials_28_0_3 & partials_28_21 |
    reducedPartials_reducedPartials_sum_475 & partials_28_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_28_0_4 = reducedPartials_reducedPartials_sum_476 ^ partials_28_22 ^
    partials_28_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_613 = reducedPartials_reducedPartials_sum_476 & partials_28_22 |
    partials_28_22 & partials_28_23 | reducedPartials_reducedPartials_sum_476 & partials_28_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_477 = reducedPartials_reducedPartials_carry_613 ^
    reducedPartials_reducedPartials_carry_612 ^ reducedPartials_reducedPartials_carry_611; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_614 = reducedPartials_reducedPartials_carry_613 &
    reducedPartials_reducedPartials_carry_612 | reducedPartials_reducedPartials_carry_612 &
    reducedPartials_reducedPartials_carry_611 | reducedPartials_reducedPartials_carry_613 &
    reducedPartials_reducedPartials_carry_611; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_478 = reducedPartials_reducedPartials_sum_477 ^
    reducedPartials_reducedPartials_29_0_3 ^ partials_29_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_615 = reducedPartials_reducedPartials_sum_477 &
    reducedPartials_reducedPartials_29_0_3 | reducedPartials_reducedPartials_29_0_3 & partials_29_22 |
    reducedPartials_reducedPartials_sum_477 & partials_29_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_29_0_4 = reducedPartials_reducedPartials_sum_478 ^ partials_29_23 ^
    partials_29_24; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_616 = reducedPartials_reducedPartials_sum_478 & partials_29_23 |
    partials_29_23 & partials_29_24 | reducedPartials_reducedPartials_sum_478 & partials_29_24; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_479 = reducedPartials_reducedPartials_carry_616 ^
    reducedPartials_reducedPartials_carry_615 ^ reducedPartials_reducedPartials_carry_614; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_617 = reducedPartials_reducedPartials_carry_616 &
    reducedPartials_reducedPartials_carry_615 | reducedPartials_reducedPartials_carry_615 &
    reducedPartials_reducedPartials_carry_614 | reducedPartials_reducedPartials_carry_616 &
    reducedPartials_reducedPartials_carry_614; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_480 = reducedPartials_reducedPartials_sum_479 ^
    reducedPartials_reducedPartials_30_0_3 ^ partials_30_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_618 = reducedPartials_reducedPartials_sum_479 &
    reducedPartials_reducedPartials_30_0_3 | reducedPartials_reducedPartials_30_0_3 & partials_30_23 |
    reducedPartials_reducedPartials_sum_479 & partials_30_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_30_0_4 = reducedPartials_reducedPartials_sum_480 ^ partials_30_24 ^
    partials_30_25; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_619 = reducedPartials_reducedPartials_sum_480 & partials_30_24 |
    partials_30_24 & partials_30_25 | reducedPartials_reducedPartials_sum_480 & partials_30_25; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_481 = reducedPartials_reducedPartials_carry_619 ^
    reducedPartials_reducedPartials_carry_618 ^ reducedPartials_reducedPartials_carry_617; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_620 = reducedPartials_reducedPartials_carry_619 &
    reducedPartials_reducedPartials_carry_618 | reducedPartials_reducedPartials_carry_618 &
    reducedPartials_reducedPartials_carry_617 | reducedPartials_reducedPartials_carry_619 &
    reducedPartials_reducedPartials_carry_617; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_482 = reducedPartials_reducedPartials_sum_481 ^
    reducedPartials_reducedPartials_31_0_3 ^ partials_31_24; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_621 = reducedPartials_reducedPartials_sum_481 &
    reducedPartials_reducedPartials_31_0_3 | reducedPartials_reducedPartials_31_0_3 & partials_31_24 |
    reducedPartials_reducedPartials_sum_481 & partials_31_24; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_31_0_4 = reducedPartials_reducedPartials_sum_482 ^ partials_31_25 ^
    partials_31_26; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_622 = reducedPartials_reducedPartials_sum_482 & partials_31_25 |
    partials_31_25 & partials_31_26 | reducedPartials_reducedPartials_sum_482 & partials_31_26; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_483 = reducedPartials_reducedPartials_carry_622 ^
    reducedPartials_reducedPartials_carry_621 ^ reducedPartials_reducedPartials_carry_620; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_623 = reducedPartials_reducedPartials_carry_622 &
    reducedPartials_reducedPartials_carry_621 | reducedPartials_reducedPartials_carry_621 &
    reducedPartials_reducedPartials_carry_620 | reducedPartials_reducedPartials_carry_622 &
    reducedPartials_reducedPartials_carry_620; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_484 = reducedPartials_reducedPartials_sum_483 ^
    reducedPartials_reducedPartials_32_0_3 ^ partials_32_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_624 = reducedPartials_reducedPartials_sum_483 &
    reducedPartials_reducedPartials_32_0_3 | reducedPartials_reducedPartials_32_0_3 & partials_32_23 |
    reducedPartials_reducedPartials_sum_483 & partials_32_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_32_0_4 = reducedPartials_reducedPartials_sum_484 ^ partials_32_24 ^
    partials_32_25; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_625 = reducedPartials_reducedPartials_sum_484 & partials_32_24 |
    partials_32_24 & partials_32_25 | reducedPartials_reducedPartials_sum_484 & partials_32_25; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_485 = reducedPartials_reducedPartials_carry_625 ^
    reducedPartials_reducedPartials_carry_624 ^ reducedPartials_reducedPartials_carry_623; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_626 = reducedPartials_reducedPartials_carry_625 &
    reducedPartials_reducedPartials_carry_624 | reducedPartials_reducedPartials_carry_624 &
    reducedPartials_reducedPartials_carry_623 | reducedPartials_reducedPartials_carry_625 &
    reducedPartials_reducedPartials_carry_623; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_486 = reducedPartials_reducedPartials_sum_485 ^
    reducedPartials_reducedPartials_33_0_3 ^ partials_33_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_627 = reducedPartials_reducedPartials_sum_485 &
    reducedPartials_reducedPartials_33_0_3 | reducedPartials_reducedPartials_33_0_3 & partials_33_22 |
    reducedPartials_reducedPartials_sum_485 & partials_33_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_33_0_4 = reducedPartials_reducedPartials_sum_486 ^ partials_33_23 ^
    partials_33_24; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_628 = reducedPartials_reducedPartials_sum_486 & partials_33_23 |
    partials_33_23 & partials_33_24 | reducedPartials_reducedPartials_sum_486 & partials_33_24; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_487 = reducedPartials_reducedPartials_carry_628 ^
    reducedPartials_reducedPartials_carry_627 ^ reducedPartials_reducedPartials_carry_626; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_629 = reducedPartials_reducedPartials_carry_628 &
    reducedPartials_reducedPartials_carry_627 | reducedPartials_reducedPartials_carry_627 &
    reducedPartials_reducedPartials_carry_626 | reducedPartials_reducedPartials_carry_628 &
    reducedPartials_reducedPartials_carry_626; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_488 = reducedPartials_reducedPartials_sum_487 ^
    reducedPartials_reducedPartials_34_0_3 ^ partials_34_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_630 = reducedPartials_reducedPartials_sum_487 &
    reducedPartials_reducedPartials_34_0_3 | reducedPartials_reducedPartials_34_0_3 & partials_34_21 |
    reducedPartials_reducedPartials_sum_487 & partials_34_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_34_0_4 = reducedPartials_reducedPartials_sum_488 ^ partials_34_22 ^
    partials_34_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_631 = reducedPartials_reducedPartials_sum_488 & partials_34_22 |
    partials_34_22 & partials_34_23 | reducedPartials_reducedPartials_sum_488 & partials_34_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_489 = reducedPartials_reducedPartials_carry_631 ^
    reducedPartials_reducedPartials_carry_630 ^ reducedPartials_reducedPartials_carry_629; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_632 = reducedPartials_reducedPartials_carry_631 &
    reducedPartials_reducedPartials_carry_630 | reducedPartials_reducedPartials_carry_630 &
    reducedPartials_reducedPartials_carry_629 | reducedPartials_reducedPartials_carry_631 &
    reducedPartials_reducedPartials_carry_629; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_490 = reducedPartials_reducedPartials_sum_489 ^
    reducedPartials_reducedPartials_35_0_3 ^ partials_35_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_633 = reducedPartials_reducedPartials_sum_489 &
    reducedPartials_reducedPartials_35_0_3 | reducedPartials_reducedPartials_35_0_3 & partials_35_20 |
    reducedPartials_reducedPartials_sum_489 & partials_35_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_35_0_4 = reducedPartials_reducedPartials_sum_490 ^ partials_35_21 ^
    partials_35_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_634 = reducedPartials_reducedPartials_sum_490 & partials_35_21 |
    partials_35_21 & partials_35_22 | reducedPartials_reducedPartials_sum_490 & partials_35_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_491 = reducedPartials_reducedPartials_carry_634 ^
    reducedPartials_reducedPartials_carry_633 ^ reducedPartials_reducedPartials_carry_632; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_635 = reducedPartials_reducedPartials_carry_634 &
    reducedPartials_reducedPartials_carry_633 | reducedPartials_reducedPartials_carry_633 &
    reducedPartials_reducedPartials_carry_632 | reducedPartials_reducedPartials_carry_634 &
    reducedPartials_reducedPartials_carry_632; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_492 = reducedPartials_reducedPartials_sum_491 ^
    reducedPartials_reducedPartials_36_0_3 ^ partials_36_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_636 = reducedPartials_reducedPartials_sum_491 &
    reducedPartials_reducedPartials_36_0_3 | reducedPartials_reducedPartials_36_0_3 & partials_36_19 |
    reducedPartials_reducedPartials_sum_491 & partials_36_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_36_0_4 = reducedPartials_reducedPartials_sum_492 ^ partials_36_20 ^
    partials_36_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_637 = reducedPartials_reducedPartials_sum_492 & partials_36_20 |
    partials_36_20 & partials_36_21 | reducedPartials_reducedPartials_sum_492 & partials_36_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_493 = reducedPartials_reducedPartials_carry_637 ^
    reducedPartials_reducedPartials_carry_636 ^ reducedPartials_reducedPartials_carry_635; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_638 = reducedPartials_reducedPartials_carry_637 &
    reducedPartials_reducedPartials_carry_636 | reducedPartials_reducedPartials_carry_636 &
    reducedPartials_reducedPartials_carry_635 | reducedPartials_reducedPartials_carry_637 &
    reducedPartials_reducedPartials_carry_635; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_494 = reducedPartials_reducedPartials_sum_493 ^
    reducedPartials_reducedPartials_37_0_2 ^ partials_37_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_639 = reducedPartials_reducedPartials_sum_493 &
    reducedPartials_reducedPartials_37_0_2 | reducedPartials_reducedPartials_37_0_2 & partials_37_18 |
    reducedPartials_reducedPartials_sum_493 & partials_37_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_37_0_3 = reducedPartials_reducedPartials_sum_494 ^ partials_37_19 ^
    partials_37_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_640 = reducedPartials_reducedPartials_sum_494 & partials_37_19 |
    partials_37_19 & partials_37_20 | reducedPartials_reducedPartials_sum_494 & partials_37_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_495 = reducedPartials_reducedPartials_carry_640 ^
    reducedPartials_reducedPartials_carry_639 ^ reducedPartials_reducedPartials_carry_638; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_641 = reducedPartials_reducedPartials_carry_640 &
    reducedPartials_reducedPartials_carry_639 | reducedPartials_reducedPartials_carry_639 &
    reducedPartials_reducedPartials_carry_638 | reducedPartials_reducedPartials_carry_640 &
    reducedPartials_reducedPartials_carry_638; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_496 = reducedPartials_reducedPartials_sum_495 ^
    reducedPartials_reducedPartials_38_0_2 ^ partials_38_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_642 = reducedPartials_reducedPartials_sum_495 &
    reducedPartials_reducedPartials_38_0_2 | reducedPartials_reducedPartials_38_0_2 & partials_38_17 |
    reducedPartials_reducedPartials_sum_495 & partials_38_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_38_0_3 = reducedPartials_reducedPartials_sum_496 ^ partials_38_18 ^
    partials_38_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_643 = reducedPartials_reducedPartials_sum_496 & partials_38_18 |
    partials_38_18 & partials_38_19 | reducedPartials_reducedPartials_sum_496 & partials_38_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_497 = reducedPartials_reducedPartials_carry_643 ^
    reducedPartials_reducedPartials_carry_642 ^ reducedPartials_reducedPartials_carry_641; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_644 = reducedPartials_reducedPartials_carry_643 &
    reducedPartials_reducedPartials_carry_642 | reducedPartials_reducedPartials_carry_642 &
    reducedPartials_reducedPartials_carry_641 | reducedPartials_reducedPartials_carry_643 &
    reducedPartials_reducedPartials_carry_641; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_498 = reducedPartials_reducedPartials_sum_497 ^
    reducedPartials_reducedPartials_39_0_2 ^ partials_39_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_645 = reducedPartials_reducedPartials_sum_497 &
    reducedPartials_reducedPartials_39_0_2 | reducedPartials_reducedPartials_39_0_2 & partials_39_16 |
    reducedPartials_reducedPartials_sum_497 & partials_39_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_39_0_3 = reducedPartials_reducedPartials_sum_498 ^ partials_39_17 ^
    partials_39_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_646 = reducedPartials_reducedPartials_sum_498 & partials_39_17 |
    partials_39_17 & partials_39_18 | reducedPartials_reducedPartials_sum_498 & partials_39_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_499 = reducedPartials_reducedPartials_carry_646 ^
    reducedPartials_reducedPartials_carry_645 ^ reducedPartials_reducedPartials_carry_644; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_647 = reducedPartials_reducedPartials_carry_646 &
    reducedPartials_reducedPartials_carry_645 | reducedPartials_reducedPartials_carry_645 &
    reducedPartials_reducedPartials_carry_644 | reducedPartials_reducedPartials_carry_646 &
    reducedPartials_reducedPartials_carry_644; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_500 = reducedPartials_reducedPartials_sum_499 ^
    reducedPartials_reducedPartials_40_0_2 ^ partials_40_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_648 = reducedPartials_reducedPartials_sum_499 &
    reducedPartials_reducedPartials_40_0_2 | reducedPartials_reducedPartials_40_0_2 & partials_40_15 |
    reducedPartials_reducedPartials_sum_499 & partials_40_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_40_0_3 = reducedPartials_reducedPartials_sum_500 ^ partials_40_16 ^
    partials_40_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_649 = reducedPartials_reducedPartials_sum_500 & partials_40_16 |
    partials_40_16 & partials_40_17 | reducedPartials_reducedPartials_sum_500 & partials_40_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_501 = reducedPartials_reducedPartials_carry_649 ^
    reducedPartials_reducedPartials_carry_648 ^ reducedPartials_reducedPartials_carry_647; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_650 = reducedPartials_reducedPartials_carry_649 &
    reducedPartials_reducedPartials_carry_648 | reducedPartials_reducedPartials_carry_648 &
    reducedPartials_reducedPartials_carry_647 | reducedPartials_reducedPartials_carry_649 &
    reducedPartials_reducedPartials_carry_647; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_502 = reducedPartials_reducedPartials_sum_501 ^
    reducedPartials_reducedPartials_41_0_2 ^ partials_41_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_651 = reducedPartials_reducedPartials_sum_501 &
    reducedPartials_reducedPartials_41_0_2 | reducedPartials_reducedPartials_41_0_2 & partials_41_14 |
    reducedPartials_reducedPartials_sum_501 & partials_41_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_41_0_3 = reducedPartials_reducedPartials_sum_502 ^ partials_41_15 ^
    partials_41_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_652 = reducedPartials_reducedPartials_sum_502 & partials_41_15 |
    partials_41_15 & partials_41_16 | reducedPartials_reducedPartials_sum_502 & partials_41_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_503 = reducedPartials_reducedPartials_carry_652 ^
    reducedPartials_reducedPartials_carry_651 ^ reducedPartials_reducedPartials_carry_650; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_653 = reducedPartials_reducedPartials_carry_652 &
    reducedPartials_reducedPartials_carry_651 | reducedPartials_reducedPartials_carry_651 &
    reducedPartials_reducedPartials_carry_650 | reducedPartials_reducedPartials_carry_652 &
    reducedPartials_reducedPartials_carry_650; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_504 = reducedPartials_reducedPartials_sum_503 ^
    reducedPartials_reducedPartials_42_0_2 ^ partials_42_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_654 = reducedPartials_reducedPartials_sum_503 &
    reducedPartials_reducedPartials_42_0_2 | reducedPartials_reducedPartials_42_0_2 & partials_42_13 |
    reducedPartials_reducedPartials_sum_503 & partials_42_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_42_0_3 = reducedPartials_reducedPartials_sum_504 ^ partials_42_14 ^
    partials_42_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_655 = reducedPartials_reducedPartials_sum_504 & partials_42_14 |
    partials_42_14 & partials_42_15 | reducedPartials_reducedPartials_sum_504 & partials_42_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_505 = reducedPartials_reducedPartials_carry_655 ^
    reducedPartials_reducedPartials_carry_654 ^ reducedPartials_reducedPartials_carry_653; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_656 = reducedPartials_reducedPartials_carry_655 &
    reducedPartials_reducedPartials_carry_654 | reducedPartials_reducedPartials_carry_654 &
    reducedPartials_reducedPartials_carry_653 | reducedPartials_reducedPartials_carry_655 &
    reducedPartials_reducedPartials_carry_653; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_506 = reducedPartials_reducedPartials_sum_505 ^
    reducedPartials_reducedPartials_43_0_2 ^ partials_43_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_657 = reducedPartials_reducedPartials_sum_505 &
    reducedPartials_reducedPartials_43_0_2 | reducedPartials_reducedPartials_43_0_2 & partials_43_12 |
    reducedPartials_reducedPartials_sum_505 & partials_43_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_43_0_3 = reducedPartials_reducedPartials_sum_506 ^ partials_43_13 ^
    partials_43_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_658 = reducedPartials_reducedPartials_sum_506 & partials_43_13 |
    partials_43_13 & partials_43_14 | reducedPartials_reducedPartials_sum_506 & partials_43_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_507 = reducedPartials_reducedPartials_carry_658 ^
    reducedPartials_reducedPartials_carry_657 ^ reducedPartials_reducedPartials_carry_656; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_659 = reducedPartials_reducedPartials_carry_658 &
    reducedPartials_reducedPartials_carry_657 | reducedPartials_reducedPartials_carry_657 &
    reducedPartials_reducedPartials_carry_656 | reducedPartials_reducedPartials_carry_658 &
    reducedPartials_reducedPartials_carry_656; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_508 = reducedPartials_reducedPartials_sum_507 ^
    reducedPartials_reducedPartials_44_0_2 ^ partials_44_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_660 = reducedPartials_reducedPartials_sum_507 &
    reducedPartials_reducedPartials_44_0_2 | reducedPartials_reducedPartials_44_0_2 & partials_44_11 |
    reducedPartials_reducedPartials_sum_507 & partials_44_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_44_0_3 = reducedPartials_reducedPartials_sum_508 ^ partials_44_12 ^
    partials_44_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_661 = reducedPartials_reducedPartials_sum_508 & partials_44_12 |
    partials_44_12 & partials_44_13 | reducedPartials_reducedPartials_sum_508 & partials_44_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_509 = reducedPartials_reducedPartials_carry_661 ^
    reducedPartials_reducedPartials_carry_660 ^ reducedPartials_reducedPartials_carry_659; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_662 = reducedPartials_reducedPartials_carry_661 &
    reducedPartials_reducedPartials_carry_660 | reducedPartials_reducedPartials_carry_660 &
    reducedPartials_reducedPartials_carry_659 | reducedPartials_reducedPartials_carry_661 &
    reducedPartials_reducedPartials_carry_659; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_510 = reducedPartials_reducedPartials_sum_509 ^
    reducedPartials_reducedPartials_45_0_2 ^ partials_45_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_663 = reducedPartials_reducedPartials_sum_509 &
    reducedPartials_reducedPartials_45_0_2 | reducedPartials_reducedPartials_45_0_2 & partials_45_10 |
    reducedPartials_reducedPartials_sum_509 & partials_45_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_45_0_3 = reducedPartials_reducedPartials_sum_510 ^ partials_45_11 ^
    partials_45_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_664 = reducedPartials_reducedPartials_sum_510 & partials_45_11 |
    partials_45_11 & partials_45_12 | reducedPartials_reducedPartials_sum_510 & partials_45_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_511 = reducedPartials_reducedPartials_carry_664 ^
    reducedPartials_reducedPartials_carry_663 ^ reducedPartials_reducedPartials_carry_662; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_665 = reducedPartials_reducedPartials_carry_664 &
    reducedPartials_reducedPartials_carry_663 | reducedPartials_reducedPartials_carry_663 &
    reducedPartials_reducedPartials_carry_662 | reducedPartials_reducedPartials_carry_664 &
    reducedPartials_reducedPartials_carry_662; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_512 = reducedPartials_reducedPartials_sum_511 ^
    reducedPartials_reducedPartials_46_0_1 ^ partials_46_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_666 = reducedPartials_reducedPartials_sum_511 &
    reducedPartials_reducedPartials_46_0_1 | reducedPartials_reducedPartials_46_0_1 & partials_46_9 |
    reducedPartials_reducedPartials_sum_511 & partials_46_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_46_0_2 = reducedPartials_reducedPartials_sum_512 ^ partials_46_10 ^
    partials_46_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_667 = reducedPartials_reducedPartials_sum_512 & partials_46_10 |
    partials_46_10 & partials_46_11 | reducedPartials_reducedPartials_sum_512 & partials_46_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_513 = reducedPartials_reducedPartials_carry_667 ^
    reducedPartials_reducedPartials_carry_666 ^ reducedPartials_reducedPartials_carry_665; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_668 = reducedPartials_reducedPartials_carry_667 &
    reducedPartials_reducedPartials_carry_666 | reducedPartials_reducedPartials_carry_666 &
    reducedPartials_reducedPartials_carry_665 | reducedPartials_reducedPartials_carry_667 &
    reducedPartials_reducedPartials_carry_665; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_514 = reducedPartials_reducedPartials_sum_513 ^
    reducedPartials_reducedPartials_47_0_1 ^ partials_47_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_669 = reducedPartials_reducedPartials_sum_513 &
    reducedPartials_reducedPartials_47_0_1 | reducedPartials_reducedPartials_47_0_1 & partials_47_8 |
    reducedPartials_reducedPartials_sum_513 & partials_47_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_47_0_2 = reducedPartials_reducedPartials_sum_514 ^ partials_47_9 ^
    partials_47_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_670 = reducedPartials_reducedPartials_sum_514 & partials_47_9 |
    partials_47_9 & partials_47_10 | reducedPartials_reducedPartials_sum_514 & partials_47_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_515 = reducedPartials_reducedPartials_carry_670 ^
    reducedPartials_reducedPartials_carry_669 ^ reducedPartials_reducedPartials_carry_668; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_671 = reducedPartials_reducedPartials_carry_670 &
    reducedPartials_reducedPartials_carry_669 | reducedPartials_reducedPartials_carry_669 &
    reducedPartials_reducedPartials_carry_668 | reducedPartials_reducedPartials_carry_670 &
    reducedPartials_reducedPartials_carry_668; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_516 = reducedPartials_reducedPartials_sum_515 ^
    reducedPartials_reducedPartials_48_0_1 ^ partials_48_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_672 = reducedPartials_reducedPartials_sum_515 &
    reducedPartials_reducedPartials_48_0_1 | reducedPartials_reducedPartials_48_0_1 & partials_48_7 |
    reducedPartials_reducedPartials_sum_515 & partials_48_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_48_0_2 = reducedPartials_reducedPartials_sum_516 ^ partials_48_8 ^ partials_48_9
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_673 = reducedPartials_reducedPartials_sum_516 & partials_48_8 |
    partials_48_8 & partials_48_9 | reducedPartials_reducedPartials_sum_516 & partials_48_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_517 = reducedPartials_reducedPartials_carry_673 ^
    reducedPartials_reducedPartials_carry_672 ^ reducedPartials_reducedPartials_carry_671; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_674 = reducedPartials_reducedPartials_carry_673 &
    reducedPartials_reducedPartials_carry_672 | reducedPartials_reducedPartials_carry_672 &
    reducedPartials_reducedPartials_carry_671 | reducedPartials_reducedPartials_carry_673 &
    reducedPartials_reducedPartials_carry_671; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_518 = reducedPartials_reducedPartials_sum_517 ^
    reducedPartials_reducedPartials_49_0_1 ^ partials_49_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_675 = reducedPartials_reducedPartials_sum_517 &
    reducedPartials_reducedPartials_49_0_1 | reducedPartials_reducedPartials_49_0_1 & partials_49_6 |
    reducedPartials_reducedPartials_sum_517 & partials_49_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_49_0_2 = reducedPartials_reducedPartials_sum_518 ^ partials_49_7 ^ partials_49_8
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_676 = reducedPartials_reducedPartials_sum_518 & partials_49_7 |
    partials_49_7 & partials_49_8 | reducedPartials_reducedPartials_sum_518 & partials_49_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_519 = reducedPartials_reducedPartials_carry_676 ^
    reducedPartials_reducedPartials_carry_675 ^ reducedPartials_reducedPartials_carry_674; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_677 = reducedPartials_reducedPartials_carry_676 &
    reducedPartials_reducedPartials_carry_675 | reducedPartials_reducedPartials_carry_675 &
    reducedPartials_reducedPartials_carry_674 | reducedPartials_reducedPartials_carry_676 &
    reducedPartials_reducedPartials_carry_674; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_520 = reducedPartials_reducedPartials_sum_519 ^
    reducedPartials_reducedPartials_50_0_1 ^ partials_50_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_678 = reducedPartials_reducedPartials_sum_519 &
    reducedPartials_reducedPartials_50_0_1 | reducedPartials_reducedPartials_50_0_1 & partials_50_5 |
    reducedPartials_reducedPartials_sum_519 & partials_50_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_50_0_2 = reducedPartials_reducedPartials_sum_520 ^ partials_50_6 ^ partials_50_7
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_679 = reducedPartials_reducedPartials_sum_520 & partials_50_6 |
    partials_50_6 & partials_50_7 | reducedPartials_reducedPartials_sum_520 & partials_50_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_521 = reducedPartials_reducedPartials_carry_679 ^
    reducedPartials_reducedPartials_carry_678 ^ reducedPartials_reducedPartials_carry_677; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_680 = reducedPartials_reducedPartials_carry_679 &
    reducedPartials_reducedPartials_carry_678 | reducedPartials_reducedPartials_carry_678 &
    reducedPartials_reducedPartials_carry_677 | reducedPartials_reducedPartials_carry_679 &
    reducedPartials_reducedPartials_carry_677; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_522 = reducedPartials_reducedPartials_sum_521 ^
    reducedPartials_reducedPartials_51_0_1 ^ partials_51_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_681 = reducedPartials_reducedPartials_sum_521 &
    reducedPartials_reducedPartials_51_0_1 | reducedPartials_reducedPartials_51_0_1 & partials_51_4 |
    reducedPartials_reducedPartials_sum_521 & partials_51_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_51_0_2 = reducedPartials_reducedPartials_sum_522 ^ partials_51_5 ^ partials_51_6
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_682 = reducedPartials_reducedPartials_sum_522 & partials_51_5 |
    partials_51_5 & partials_51_6 | reducedPartials_reducedPartials_sum_522 & partials_51_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_523 = reducedPartials_reducedPartials_carry_682 ^
    reducedPartials_reducedPartials_carry_681 ^ reducedPartials_reducedPartials_carry_680; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_683 = reducedPartials_reducedPartials_carry_682 &
    reducedPartials_reducedPartials_carry_681 | reducedPartials_reducedPartials_carry_681 &
    reducedPartials_reducedPartials_carry_680 | reducedPartials_reducedPartials_carry_682 &
    reducedPartials_reducedPartials_carry_680; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_524 = reducedPartials_reducedPartials_sum_523 ^
    reducedPartials_reducedPartials_52_0 ^ partials_52_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_684 = reducedPartials_reducedPartials_sum_523 &
    reducedPartials_reducedPartials_52_0 | reducedPartials_reducedPartials_52_0 & partials_52_3 |
    reducedPartials_reducedPartials_sum_523 & partials_52_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_52_0_1 = reducedPartials_reducedPartials_sum_524 ^ partials_52_4 ^ partials_52_5
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_685 = reducedPartials_reducedPartials_sum_524 & partials_52_4 |
    partials_52_4 & partials_52_5 | reducedPartials_reducedPartials_sum_524 & partials_52_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_525 = reducedPartials_reducedPartials_carry_685 ^
    reducedPartials_reducedPartials_carry_684 ^ reducedPartials_reducedPartials_carry_683; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_686 = reducedPartials_reducedPartials_carry_685 &
    reducedPartials_reducedPartials_carry_684 | reducedPartials_reducedPartials_carry_684 &
    reducedPartials_reducedPartials_carry_683 | reducedPartials_reducedPartials_carry_685 &
    reducedPartials_reducedPartials_carry_683; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_526 = reducedPartials_reducedPartials_sum_525 ^
    reducedPartials_reducedPartials_53_0 ^ partials_53_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_687 = reducedPartials_reducedPartials_sum_525 &
    reducedPartials_reducedPartials_53_0 | reducedPartials_reducedPartials_53_0 & partials_53_2 |
    reducedPartials_reducedPartials_sum_525 & partials_53_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_53_0_1 = reducedPartials_reducedPartials_sum_526 ^ partials_53_3 ^ partials_53_4
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_688 = reducedPartials_reducedPartials_sum_526 & partials_53_3 |
    partials_53_3 & partials_53_4 | reducedPartials_reducedPartials_sum_526 & partials_53_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_527 = reducedPartials_reducedPartials_carry_688 ^
    reducedPartials_reducedPartials_carry_687 ^ reducedPartials_reducedPartials_carry_686; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_689 = reducedPartials_reducedPartials_carry_688 &
    reducedPartials_reducedPartials_carry_687 | reducedPartials_reducedPartials_carry_687 &
    reducedPartials_reducedPartials_carry_686 | reducedPartials_reducedPartials_carry_688 &
    reducedPartials_reducedPartials_carry_686; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_528 = reducedPartials_reducedPartials_sum_527 ^
    reducedPartials_reducedPartials_54_0 ^ partials_54_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_690 = reducedPartials_reducedPartials_sum_527 &
    reducedPartials_reducedPartials_54_0 | reducedPartials_reducedPartials_54_0 & partials_54_1 |
    reducedPartials_reducedPartials_sum_527 & partials_54_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_54_0_1 = reducedPartials_reducedPartials_sum_528 ^ partials_54_2 ^ partials_54_3
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_691 = reducedPartials_reducedPartials_sum_528 & partials_54_2 |
    partials_54_2 & partials_54_3 | reducedPartials_reducedPartials_sum_528 & partials_54_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_529 = reducedPartials_reducedPartials_carry_691 ^
    reducedPartials_reducedPartials_carry_690 ^ reducedPartials_reducedPartials_carry_689; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_692 = reducedPartials_reducedPartials_carry_691 &
    reducedPartials_reducedPartials_carry_690 | reducedPartials_reducedPartials_carry_690 &
    reducedPartials_reducedPartials_carry_689 | reducedPartials_reducedPartials_carry_691 &
    reducedPartials_reducedPartials_carry_689; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_530 = reducedPartials_reducedPartials_sum_529 ^
    reducedPartials_reducedPartials_55_0 ^ partials_55_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_693 = reducedPartials_reducedPartials_sum_529 &
    reducedPartials_reducedPartials_55_0 | reducedPartials_reducedPartials_55_0 & partials_55_0 |
    reducedPartials_reducedPartials_sum_529 & partials_55_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_55_0_1 = reducedPartials_reducedPartials_sum_530 ^ partials_55_1 ^ partials_55_2
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_694 = reducedPartials_reducedPartials_sum_530 & partials_55_1 |
    partials_55_1 & partials_55_2 | reducedPartials_reducedPartials_sum_530 & partials_55_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_531 = reducedPartials_reducedPartials_carry_694 ^
    reducedPartials_reducedPartials_carry_693 ^ reducedPartials_reducedPartials_carry_692; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_695 = reducedPartials_reducedPartials_carry_694 &
    reducedPartials_reducedPartials_carry_693 | reducedPartials_reducedPartials_carry_693 &
    reducedPartials_reducedPartials_carry_692 | reducedPartials_reducedPartials_carry_694 &
    reducedPartials_reducedPartials_carry_692; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_56_0 = reducedPartials_reducedPartials_sum_531 ^ partials_56_0 ^ partials_56_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_696 = reducedPartials_reducedPartials_sum_531 & partials_56_0 |
    partials_56_0 & partials_56_1 | reducedPartials_reducedPartials_sum_531 & partials_56_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_57_0 = reducedPartials_reducedPartials_carry_696 ^
    reducedPartials_reducedPartials_carry_695 ^ partials_57_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_58_0 = reducedPartials_reducedPartials_carry_696 &
    reducedPartials_reducedPartials_carry_695 | reducedPartials_reducedPartials_carry_695 & partials_57_0 |
    reducedPartials_reducedPartials_carry_696 & partials_57_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_4_0 = partials_4_0 ^ partials_4_1; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_697 = partials_4_0 & partials_4_1; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_532 = reducedPartials_reducedPartials_carry_697 ^ partials_5_0 ^
    partials_5_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_698 = reducedPartials_reducedPartials_carry_697 & partials_5_0 |
    partials_5_0 & partials_5_1 | reducedPartials_reducedPartials_carry_697 & partials_5_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_5_0 = reducedPartials_reducedPartials_sum_532 ^ partials_5_2; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_699 = reducedPartials_reducedPartials_sum_532 & partials_5_2; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_sum_533 = reducedPartials_reducedPartials_carry_699 ^
    reducedPartials_reducedPartials_carry_698 ^ reducedPartials_reducedPartials_6_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_700 = reducedPartials_reducedPartials_carry_699 &
    reducedPartials_reducedPartials_carry_698 | reducedPartials_reducedPartials_carry_698 &
    reducedPartials_reducedPartials_6_0 | reducedPartials_reducedPartials_carry_699 &
    reducedPartials_reducedPartials_6_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_6_0_1 = reducedPartials_reducedPartials_sum_533 ^ partials_6_2 ^ partials_6_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_701 = reducedPartials_reducedPartials_sum_533 & partials_6_2 |
    partials_6_2 & partials_6_3 | reducedPartials_reducedPartials_sum_533 & partials_6_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_534 = reducedPartials_reducedPartials_carry_701 ^
    reducedPartials_reducedPartials_carry_700 ^ reducedPartials_reducedPartials_7_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_702 = reducedPartials_reducedPartials_carry_701 &
    reducedPartials_reducedPartials_carry_700 | reducedPartials_reducedPartials_carry_700 &
    reducedPartials_reducedPartials_7_0 | reducedPartials_reducedPartials_carry_701 &
    reducedPartials_reducedPartials_7_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_7_0_1 = reducedPartials_reducedPartials_sum_534 ^ partials_7_3 ^ partials_7_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_703 = reducedPartials_reducedPartials_sum_534 & partials_7_3 |
    partials_7_3 & partials_7_4 | reducedPartials_reducedPartials_sum_534 & partials_7_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_535 = reducedPartials_reducedPartials_carry_703 ^
    reducedPartials_reducedPartials_carry_702 ^ reducedPartials_reducedPartials_8_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_704 = reducedPartials_reducedPartials_carry_703 &
    reducedPartials_reducedPartials_carry_702 | reducedPartials_reducedPartials_carry_702 &
    reducedPartials_reducedPartials_8_0 | reducedPartials_reducedPartials_carry_703 &
    reducedPartials_reducedPartials_8_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_8_0_1 = reducedPartials_reducedPartials_sum_535 ^ partials_8_4 ^ partials_8_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_705 = reducedPartials_reducedPartials_sum_535 & partials_8_4 |
    partials_8_4 & partials_8_5 | reducedPartials_reducedPartials_sum_535 & partials_8_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_536 = reducedPartials_reducedPartials_carry_705 ^
    reducedPartials_reducedPartials_carry_704 ^ reducedPartials_reducedPartials_9_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_706 = reducedPartials_reducedPartials_carry_705 &
    reducedPartials_reducedPartials_carry_704 | reducedPartials_reducedPartials_carry_704 &
    reducedPartials_reducedPartials_9_0_1 | reducedPartials_reducedPartials_carry_705 &
    reducedPartials_reducedPartials_9_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_9_0_2 = reducedPartials_reducedPartials_sum_536 ^ partials_9_5 ^ partials_9_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_707 = reducedPartials_reducedPartials_sum_536 & partials_9_5 |
    partials_9_5 & partials_9_6 | reducedPartials_reducedPartials_sum_536 & partials_9_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_537 = reducedPartials_reducedPartials_carry_707 ^
    reducedPartials_reducedPartials_carry_706 ^ reducedPartials_reducedPartials_10_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_708 = reducedPartials_reducedPartials_carry_707 &
    reducedPartials_reducedPartials_carry_706 | reducedPartials_reducedPartials_carry_706 &
    reducedPartials_reducedPartials_10_0_1 | reducedPartials_reducedPartials_carry_707 &
    reducedPartials_reducedPartials_10_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_10_0_2 = reducedPartials_reducedPartials_sum_537 ^ partials_10_6 ^ partials_10_7
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_709 = reducedPartials_reducedPartials_sum_537 & partials_10_6 |
    partials_10_6 & partials_10_7 | reducedPartials_reducedPartials_sum_537 & partials_10_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_538 = reducedPartials_reducedPartials_carry_709 ^
    reducedPartials_reducedPartials_carry_708 ^ reducedPartials_reducedPartials_11_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_710 = reducedPartials_reducedPartials_carry_709 &
    reducedPartials_reducedPartials_carry_708 | reducedPartials_reducedPartials_carry_708 &
    reducedPartials_reducedPartials_11_0_1 | reducedPartials_reducedPartials_carry_709 &
    reducedPartials_reducedPartials_11_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_11_0_2 = reducedPartials_reducedPartials_sum_538 ^ partials_11_7 ^ partials_11_8
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_711 = reducedPartials_reducedPartials_sum_538 & partials_11_7 |
    partials_11_7 & partials_11_8 | reducedPartials_reducedPartials_sum_538 & partials_11_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_539 = reducedPartials_reducedPartials_carry_711 ^
    reducedPartials_reducedPartials_carry_710 ^ reducedPartials_reducedPartials_12_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_712 = reducedPartials_reducedPartials_carry_711 &
    reducedPartials_reducedPartials_carry_710 | reducedPartials_reducedPartials_carry_710 &
    reducedPartials_reducedPartials_12_0_1 | reducedPartials_reducedPartials_carry_711 &
    reducedPartials_reducedPartials_12_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_12_0_2 = reducedPartials_reducedPartials_sum_539 ^ partials_12_8 ^ partials_12_9
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_713 = reducedPartials_reducedPartials_sum_539 & partials_12_8 |
    partials_12_8 & partials_12_9 | reducedPartials_reducedPartials_sum_539 & partials_12_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_540 = reducedPartials_reducedPartials_carry_713 ^
    reducedPartials_reducedPartials_carry_712 ^ reducedPartials_reducedPartials_13_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_714 = reducedPartials_reducedPartials_carry_713 &
    reducedPartials_reducedPartials_carry_712 | reducedPartials_reducedPartials_carry_712 &
    reducedPartials_reducedPartials_13_0_2 | reducedPartials_reducedPartials_carry_713 &
    reducedPartials_reducedPartials_13_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_13_0_3 = reducedPartials_reducedPartials_sum_540 ^ partials_13_9 ^
    partials_13_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_715 = reducedPartials_reducedPartials_sum_540 & partials_13_9 |
    partials_13_9 & partials_13_10 | reducedPartials_reducedPartials_sum_540 & partials_13_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_541 = reducedPartials_reducedPartials_carry_715 ^
    reducedPartials_reducedPartials_carry_714 ^ reducedPartials_reducedPartials_14_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_716 = reducedPartials_reducedPartials_carry_715 &
    reducedPartials_reducedPartials_carry_714 | reducedPartials_reducedPartials_carry_714 &
    reducedPartials_reducedPartials_14_0_2 | reducedPartials_reducedPartials_carry_715 &
    reducedPartials_reducedPartials_14_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_14_0_3 = reducedPartials_reducedPartials_sum_541 ^ partials_14_10 ^
    partials_14_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_717 = reducedPartials_reducedPartials_sum_541 & partials_14_10 |
    partials_14_10 & partials_14_11 | reducedPartials_reducedPartials_sum_541 & partials_14_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_542 = reducedPartials_reducedPartials_carry_717 ^
    reducedPartials_reducedPartials_carry_716 ^ reducedPartials_reducedPartials_15_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_718 = reducedPartials_reducedPartials_carry_717 &
    reducedPartials_reducedPartials_carry_716 | reducedPartials_reducedPartials_carry_716 &
    reducedPartials_reducedPartials_15_0_2 | reducedPartials_reducedPartials_carry_717 &
    reducedPartials_reducedPartials_15_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_15_0_3 = reducedPartials_reducedPartials_sum_542 ^ partials_15_11 ^
    partials_15_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_719 = reducedPartials_reducedPartials_sum_542 & partials_15_11 |
    partials_15_11 & partials_15_12 | reducedPartials_reducedPartials_sum_542 & partials_15_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_543 = reducedPartials_reducedPartials_carry_719 ^
    reducedPartials_reducedPartials_carry_718 ^ reducedPartials_reducedPartials_16_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_720 = reducedPartials_reducedPartials_carry_719 &
    reducedPartials_reducedPartials_carry_718 | reducedPartials_reducedPartials_carry_718 &
    reducedPartials_reducedPartials_16_0_2 | reducedPartials_reducedPartials_carry_719 &
    reducedPartials_reducedPartials_16_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_16_0_3 = reducedPartials_reducedPartials_sum_543 ^ partials_16_12 ^
    partials_16_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_721 = reducedPartials_reducedPartials_sum_543 & partials_16_12 |
    partials_16_12 & partials_16_13 | reducedPartials_reducedPartials_sum_543 & partials_16_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_544 = reducedPartials_reducedPartials_carry_721 ^
    reducedPartials_reducedPartials_carry_720 ^ reducedPartials_reducedPartials_17_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_722 = reducedPartials_reducedPartials_carry_721 &
    reducedPartials_reducedPartials_carry_720 | reducedPartials_reducedPartials_carry_720 &
    reducedPartials_reducedPartials_17_0_2 | reducedPartials_reducedPartials_carry_721 &
    reducedPartials_reducedPartials_17_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_17_0_3 = reducedPartials_reducedPartials_sum_544 ^ partials_17_13 ^
    partials_17_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_723 = reducedPartials_reducedPartials_sum_544 & partials_17_13 |
    partials_17_13 & partials_17_14 | reducedPartials_reducedPartials_sum_544 & partials_17_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_545 = reducedPartials_reducedPartials_carry_723 ^
    reducedPartials_reducedPartials_carry_722 ^ reducedPartials_reducedPartials_18_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_724 = reducedPartials_reducedPartials_carry_723 &
    reducedPartials_reducedPartials_carry_722 | reducedPartials_reducedPartials_carry_722 &
    reducedPartials_reducedPartials_18_0_2 | reducedPartials_reducedPartials_carry_723 &
    reducedPartials_reducedPartials_18_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_18_0_3 = reducedPartials_reducedPartials_sum_545 ^ partials_18_14 ^
    partials_18_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_725 = reducedPartials_reducedPartials_sum_545 & partials_18_14 |
    partials_18_14 & partials_18_15 | reducedPartials_reducedPartials_sum_545 & partials_18_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_546 = reducedPartials_reducedPartials_carry_725 ^
    reducedPartials_reducedPartials_carry_724 ^ reducedPartials_reducedPartials_19_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_726 = reducedPartials_reducedPartials_carry_725 &
    reducedPartials_reducedPartials_carry_724 | reducedPartials_reducedPartials_carry_724 &
    reducedPartials_reducedPartials_19_0_3 | reducedPartials_reducedPartials_carry_725 &
    reducedPartials_reducedPartials_19_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_19_0_4 = reducedPartials_reducedPartials_sum_546 ^ partials_19_15 ^
    partials_19_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_727 = reducedPartials_reducedPartials_sum_546 & partials_19_15 |
    partials_19_15 & partials_19_16 | reducedPartials_reducedPartials_sum_546 & partials_19_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_547 = reducedPartials_reducedPartials_carry_727 ^
    reducedPartials_reducedPartials_carry_726 ^ reducedPartials_reducedPartials_20_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_728 = reducedPartials_reducedPartials_carry_727 &
    reducedPartials_reducedPartials_carry_726 | reducedPartials_reducedPartials_carry_726 &
    reducedPartials_reducedPartials_20_0_3 | reducedPartials_reducedPartials_carry_727 &
    reducedPartials_reducedPartials_20_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_20_0_4 = reducedPartials_reducedPartials_sum_547 ^ partials_20_16 ^
    partials_20_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_729 = reducedPartials_reducedPartials_sum_547 & partials_20_16 |
    partials_20_16 & partials_20_17 | reducedPartials_reducedPartials_sum_547 & partials_20_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_548 = reducedPartials_reducedPartials_carry_729 ^
    reducedPartials_reducedPartials_carry_728 ^ reducedPartials_reducedPartials_21_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_730 = reducedPartials_reducedPartials_carry_729 &
    reducedPartials_reducedPartials_carry_728 | reducedPartials_reducedPartials_carry_728 &
    reducedPartials_reducedPartials_21_0_3 | reducedPartials_reducedPartials_carry_729 &
    reducedPartials_reducedPartials_21_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_21_0_4 = reducedPartials_reducedPartials_sum_548 ^ partials_21_17 ^
    partials_21_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_731 = reducedPartials_reducedPartials_sum_548 & partials_21_17 |
    partials_21_17 & partials_21_18 | reducedPartials_reducedPartials_sum_548 & partials_21_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_549 = reducedPartials_reducedPartials_carry_731 ^
    reducedPartials_reducedPartials_carry_730 ^ reducedPartials_reducedPartials_22_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_732 = reducedPartials_reducedPartials_carry_731 &
    reducedPartials_reducedPartials_carry_730 | reducedPartials_reducedPartials_carry_730 &
    reducedPartials_reducedPartials_22_0_3 | reducedPartials_reducedPartials_carry_731 &
    reducedPartials_reducedPartials_22_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_22_0_4 = reducedPartials_reducedPartials_sum_549 ^ partials_22_18 ^
    partials_22_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_733 = reducedPartials_reducedPartials_sum_549 & partials_22_18 |
    partials_22_18 & partials_22_19 | reducedPartials_reducedPartials_sum_549 & partials_22_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_550 = reducedPartials_reducedPartials_carry_733 ^
    reducedPartials_reducedPartials_carry_732 ^ reducedPartials_reducedPartials_23_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_734 = reducedPartials_reducedPartials_carry_733 &
    reducedPartials_reducedPartials_carry_732 | reducedPartials_reducedPartials_carry_732 &
    reducedPartials_reducedPartials_23_0_3 | reducedPartials_reducedPartials_carry_733 &
    reducedPartials_reducedPartials_23_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_23_0_4 = reducedPartials_reducedPartials_sum_550 ^ partials_23_19 ^
    partials_23_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_735 = reducedPartials_reducedPartials_sum_550 & partials_23_19 |
    partials_23_19 & partials_23_20 | reducedPartials_reducedPartials_sum_550 & partials_23_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_551 = reducedPartials_reducedPartials_carry_735 ^
    reducedPartials_reducedPartials_carry_734 ^ reducedPartials_reducedPartials_24_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_736 = reducedPartials_reducedPartials_carry_735 &
    reducedPartials_reducedPartials_carry_734 | reducedPartials_reducedPartials_carry_734 &
    reducedPartials_reducedPartials_24_0_3 | reducedPartials_reducedPartials_carry_735 &
    reducedPartials_reducedPartials_24_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_24_0_4 = reducedPartials_reducedPartials_sum_551 ^ partials_24_20 ^
    partials_24_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_737 = reducedPartials_reducedPartials_sum_551 & partials_24_20 |
    partials_24_20 & partials_24_21 | reducedPartials_reducedPartials_sum_551 & partials_24_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_552 = reducedPartials_reducedPartials_carry_737 ^
    reducedPartials_reducedPartials_carry_736 ^ reducedPartials_reducedPartials_25_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_738 = reducedPartials_reducedPartials_carry_737 &
    reducedPartials_reducedPartials_carry_736 | reducedPartials_reducedPartials_carry_736 &
    reducedPartials_reducedPartials_25_0_3 | reducedPartials_reducedPartials_carry_737 &
    reducedPartials_reducedPartials_25_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_25_0_4 = reducedPartials_reducedPartials_sum_552 ^ partials_25_21 ^
    partials_25_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_739 = reducedPartials_reducedPartials_sum_552 & partials_25_21 |
    partials_25_21 & partials_25_22 | reducedPartials_reducedPartials_sum_552 & partials_25_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_553 = reducedPartials_reducedPartials_carry_739 ^
    reducedPartials_reducedPartials_carry_738 ^ reducedPartials_reducedPartials_26_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_740 = reducedPartials_reducedPartials_carry_739 &
    reducedPartials_reducedPartials_carry_738 | reducedPartials_reducedPartials_carry_738 &
    reducedPartials_reducedPartials_26_0_3 | reducedPartials_reducedPartials_carry_739 &
    reducedPartials_reducedPartials_26_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_26_0_4 = reducedPartials_reducedPartials_sum_553 ^ partials_26_22 ^
    partials_26_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_741 = reducedPartials_reducedPartials_sum_553 & partials_26_22 |
    partials_26_22 & partials_26_23 | reducedPartials_reducedPartials_sum_553 & partials_26_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_554 = reducedPartials_reducedPartials_carry_741 ^
    reducedPartials_reducedPartials_carry_740 ^ reducedPartials_reducedPartials_27_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_742 = reducedPartials_reducedPartials_carry_741 &
    reducedPartials_reducedPartials_carry_740 | reducedPartials_reducedPartials_carry_740 &
    reducedPartials_reducedPartials_27_0_3 | reducedPartials_reducedPartials_carry_741 &
    reducedPartials_reducedPartials_27_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_27_0_4 = reducedPartials_reducedPartials_sum_554 ^ partials_27_23 ^
    partials_27_24; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_743 = reducedPartials_reducedPartials_sum_554 & partials_27_23 |
    partials_27_23 & partials_27_24 | reducedPartials_reducedPartials_sum_554 & partials_27_24; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_555 = reducedPartials_reducedPartials_carry_743 ^
    reducedPartials_reducedPartials_carry_742 ^ reducedPartials_reducedPartials_28_0_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_744 = reducedPartials_reducedPartials_carry_743 &
    reducedPartials_reducedPartials_carry_742 | reducedPartials_reducedPartials_carry_742 &
    reducedPartials_reducedPartials_28_0_4 | reducedPartials_reducedPartials_carry_743 &
    reducedPartials_reducedPartials_28_0_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_28_0_5 = reducedPartials_reducedPartials_sum_555 ^ partials_28_24 ^
    partials_28_25; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_745 = reducedPartials_reducedPartials_sum_555 & partials_28_24 |
    partials_28_24 & partials_28_25 | reducedPartials_reducedPartials_sum_555 & partials_28_25; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_556 = reducedPartials_reducedPartials_carry_745 ^
    reducedPartials_reducedPartials_carry_744 ^ reducedPartials_reducedPartials_29_0_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_746 = reducedPartials_reducedPartials_carry_745 &
    reducedPartials_reducedPartials_carry_744 | reducedPartials_reducedPartials_carry_744 &
    reducedPartials_reducedPartials_29_0_4 | reducedPartials_reducedPartials_carry_745 &
    reducedPartials_reducedPartials_29_0_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_29_0_5 = reducedPartials_reducedPartials_sum_556 ^ partials_29_25 ^
    partials_29_26; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_747 = reducedPartials_reducedPartials_sum_556 & partials_29_25 |
    partials_29_25 & partials_29_26 | reducedPartials_reducedPartials_sum_556 & partials_29_26; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_557 = reducedPartials_reducedPartials_carry_747 ^
    reducedPartials_reducedPartials_carry_746 ^ reducedPartials_reducedPartials_30_0_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_748 = reducedPartials_reducedPartials_carry_747 &
    reducedPartials_reducedPartials_carry_746 | reducedPartials_reducedPartials_carry_746 &
    reducedPartials_reducedPartials_30_0_4 | reducedPartials_reducedPartials_carry_747 &
    reducedPartials_reducedPartials_30_0_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_30_0_5 = reducedPartials_reducedPartials_sum_557 ^ partials_30_26 ^
    partials_30_27; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_749 = reducedPartials_reducedPartials_sum_557 & partials_30_26 |
    partials_30_26 & partials_30_27 | reducedPartials_reducedPartials_sum_557 & partials_30_27; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_558 = reducedPartials_reducedPartials_carry_749 ^
    reducedPartials_reducedPartials_carry_748 ^ reducedPartials_reducedPartials_31_0_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_750 = reducedPartials_reducedPartials_carry_749 &
    reducedPartials_reducedPartials_carry_748 | reducedPartials_reducedPartials_carry_748 &
    reducedPartials_reducedPartials_31_0_4 | reducedPartials_reducedPartials_carry_749 &
    reducedPartials_reducedPartials_31_0_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_31_0_5 = reducedPartials_reducedPartials_sum_558 ^ partials_31_27 ^
    partials_31_28; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_751 = reducedPartials_reducedPartials_sum_558 & partials_31_27 |
    partials_31_27 & partials_31_28 | reducedPartials_reducedPartials_sum_558 & partials_31_28; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_559 = reducedPartials_reducedPartials_carry_751 ^
    reducedPartials_reducedPartials_carry_750 ^ reducedPartials_reducedPartials_32_0_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_752 = reducedPartials_reducedPartials_carry_751 &
    reducedPartials_reducedPartials_carry_750 | reducedPartials_reducedPartials_carry_750 &
    reducedPartials_reducedPartials_32_0_4 | reducedPartials_reducedPartials_carry_751 &
    reducedPartials_reducedPartials_32_0_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_32_0_5 = reducedPartials_reducedPartials_sum_559 ^ partials_32_26 ^
    partials_32_27; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_753 = reducedPartials_reducedPartials_sum_559 & partials_32_26 |
    partials_32_26 & partials_32_27 | reducedPartials_reducedPartials_sum_559 & partials_32_27; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_560 = reducedPartials_reducedPartials_carry_753 ^
    reducedPartials_reducedPartials_carry_752 ^ reducedPartials_reducedPartials_33_0_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_754 = reducedPartials_reducedPartials_carry_753 &
    reducedPartials_reducedPartials_carry_752 | reducedPartials_reducedPartials_carry_752 &
    reducedPartials_reducedPartials_33_0_4 | reducedPartials_reducedPartials_carry_753 &
    reducedPartials_reducedPartials_33_0_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_33_0_5 = reducedPartials_reducedPartials_sum_560 ^ partials_33_25 ^
    partials_33_26; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_755 = reducedPartials_reducedPartials_sum_560 & partials_33_25 |
    partials_33_25 & partials_33_26 | reducedPartials_reducedPartials_sum_560 & partials_33_26; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_561 = reducedPartials_reducedPartials_carry_755 ^
    reducedPartials_reducedPartials_carry_754 ^ reducedPartials_reducedPartials_34_0_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_756 = reducedPartials_reducedPartials_carry_755 &
    reducedPartials_reducedPartials_carry_754 | reducedPartials_reducedPartials_carry_754 &
    reducedPartials_reducedPartials_34_0_4 | reducedPartials_reducedPartials_carry_755 &
    reducedPartials_reducedPartials_34_0_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_34_0_5 = reducedPartials_reducedPartials_sum_561 ^ partials_34_24 ^
    partials_34_25; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_757 = reducedPartials_reducedPartials_sum_561 & partials_34_24 |
    partials_34_24 & partials_34_25 | reducedPartials_reducedPartials_sum_561 & partials_34_25; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_562 = reducedPartials_reducedPartials_carry_757 ^
    reducedPartials_reducedPartials_carry_756 ^ reducedPartials_reducedPartials_35_0_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_758 = reducedPartials_reducedPartials_carry_757 &
    reducedPartials_reducedPartials_carry_756 | reducedPartials_reducedPartials_carry_756 &
    reducedPartials_reducedPartials_35_0_4 | reducedPartials_reducedPartials_carry_757 &
    reducedPartials_reducedPartials_35_0_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_35_0_5 = reducedPartials_reducedPartials_sum_562 ^ partials_35_23 ^
    partials_35_24; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_759 = reducedPartials_reducedPartials_sum_562 & partials_35_23 |
    partials_35_23 & partials_35_24 | reducedPartials_reducedPartials_sum_562 & partials_35_24; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_563 = reducedPartials_reducedPartials_carry_759 ^
    reducedPartials_reducedPartials_carry_758 ^ reducedPartials_reducedPartials_36_0_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_760 = reducedPartials_reducedPartials_carry_759 &
    reducedPartials_reducedPartials_carry_758 | reducedPartials_reducedPartials_carry_758 &
    reducedPartials_reducedPartials_36_0_4 | reducedPartials_reducedPartials_carry_759 &
    reducedPartials_reducedPartials_36_0_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_36_0_5 = reducedPartials_reducedPartials_sum_563 ^ partials_36_22 ^
    partials_36_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_761 = reducedPartials_reducedPartials_sum_563 & partials_36_22 |
    partials_36_22 & partials_36_23 | reducedPartials_reducedPartials_sum_563 & partials_36_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_564 = reducedPartials_reducedPartials_carry_761 ^
    reducedPartials_reducedPartials_carry_760 ^ reducedPartials_reducedPartials_37_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_762 = reducedPartials_reducedPartials_carry_761 &
    reducedPartials_reducedPartials_carry_760 | reducedPartials_reducedPartials_carry_760 &
    reducedPartials_reducedPartials_37_0_3 | reducedPartials_reducedPartials_carry_761 &
    reducedPartials_reducedPartials_37_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_37_0_4 = reducedPartials_reducedPartials_sum_564 ^ partials_37_21 ^
    partials_37_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_763 = reducedPartials_reducedPartials_sum_564 & partials_37_21 |
    partials_37_21 & partials_37_22 | reducedPartials_reducedPartials_sum_564 & partials_37_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_565 = reducedPartials_reducedPartials_carry_763 ^
    reducedPartials_reducedPartials_carry_762 ^ reducedPartials_reducedPartials_38_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_764 = reducedPartials_reducedPartials_carry_763 &
    reducedPartials_reducedPartials_carry_762 | reducedPartials_reducedPartials_carry_762 &
    reducedPartials_reducedPartials_38_0_3 | reducedPartials_reducedPartials_carry_763 &
    reducedPartials_reducedPartials_38_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_38_0_4 = reducedPartials_reducedPartials_sum_565 ^ partials_38_20 ^
    partials_38_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_765 = reducedPartials_reducedPartials_sum_565 & partials_38_20 |
    partials_38_20 & partials_38_21 | reducedPartials_reducedPartials_sum_565 & partials_38_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_566 = reducedPartials_reducedPartials_carry_765 ^
    reducedPartials_reducedPartials_carry_764 ^ reducedPartials_reducedPartials_39_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_766 = reducedPartials_reducedPartials_carry_765 &
    reducedPartials_reducedPartials_carry_764 | reducedPartials_reducedPartials_carry_764 &
    reducedPartials_reducedPartials_39_0_3 | reducedPartials_reducedPartials_carry_765 &
    reducedPartials_reducedPartials_39_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_39_0_4 = reducedPartials_reducedPartials_sum_566 ^ partials_39_19 ^
    partials_39_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_767 = reducedPartials_reducedPartials_sum_566 & partials_39_19 |
    partials_39_19 & partials_39_20 | reducedPartials_reducedPartials_sum_566 & partials_39_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_567 = reducedPartials_reducedPartials_carry_767 ^
    reducedPartials_reducedPartials_carry_766 ^ reducedPartials_reducedPartials_40_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_768 = reducedPartials_reducedPartials_carry_767 &
    reducedPartials_reducedPartials_carry_766 | reducedPartials_reducedPartials_carry_766 &
    reducedPartials_reducedPartials_40_0_3 | reducedPartials_reducedPartials_carry_767 &
    reducedPartials_reducedPartials_40_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_40_0_4 = reducedPartials_reducedPartials_sum_567 ^ partials_40_18 ^
    partials_40_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_769 = reducedPartials_reducedPartials_sum_567 & partials_40_18 |
    partials_40_18 & partials_40_19 | reducedPartials_reducedPartials_sum_567 & partials_40_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_568 = reducedPartials_reducedPartials_carry_769 ^
    reducedPartials_reducedPartials_carry_768 ^ reducedPartials_reducedPartials_41_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_770 = reducedPartials_reducedPartials_carry_769 &
    reducedPartials_reducedPartials_carry_768 | reducedPartials_reducedPartials_carry_768 &
    reducedPartials_reducedPartials_41_0_3 | reducedPartials_reducedPartials_carry_769 &
    reducedPartials_reducedPartials_41_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_41_0_4 = reducedPartials_reducedPartials_sum_568 ^ partials_41_17 ^
    partials_41_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_771 = reducedPartials_reducedPartials_sum_568 & partials_41_17 |
    partials_41_17 & partials_41_18 | reducedPartials_reducedPartials_sum_568 & partials_41_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_569 = reducedPartials_reducedPartials_carry_771 ^
    reducedPartials_reducedPartials_carry_770 ^ reducedPartials_reducedPartials_42_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_772 = reducedPartials_reducedPartials_carry_771 &
    reducedPartials_reducedPartials_carry_770 | reducedPartials_reducedPartials_carry_770 &
    reducedPartials_reducedPartials_42_0_3 | reducedPartials_reducedPartials_carry_771 &
    reducedPartials_reducedPartials_42_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_42_0_4 = reducedPartials_reducedPartials_sum_569 ^ partials_42_16 ^
    partials_42_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_773 = reducedPartials_reducedPartials_sum_569 & partials_42_16 |
    partials_42_16 & partials_42_17 | reducedPartials_reducedPartials_sum_569 & partials_42_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_570 = reducedPartials_reducedPartials_carry_773 ^
    reducedPartials_reducedPartials_carry_772 ^ reducedPartials_reducedPartials_43_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_774 = reducedPartials_reducedPartials_carry_773 &
    reducedPartials_reducedPartials_carry_772 | reducedPartials_reducedPartials_carry_772 &
    reducedPartials_reducedPartials_43_0_3 | reducedPartials_reducedPartials_carry_773 &
    reducedPartials_reducedPartials_43_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_43_0_4 = reducedPartials_reducedPartials_sum_570 ^ partials_43_15 ^
    partials_43_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_775 = reducedPartials_reducedPartials_sum_570 & partials_43_15 |
    partials_43_15 & partials_43_16 | reducedPartials_reducedPartials_sum_570 & partials_43_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_571 = reducedPartials_reducedPartials_carry_775 ^
    reducedPartials_reducedPartials_carry_774 ^ reducedPartials_reducedPartials_44_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_776 = reducedPartials_reducedPartials_carry_775 &
    reducedPartials_reducedPartials_carry_774 | reducedPartials_reducedPartials_carry_774 &
    reducedPartials_reducedPartials_44_0_3 | reducedPartials_reducedPartials_carry_775 &
    reducedPartials_reducedPartials_44_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_44_0_4 = reducedPartials_reducedPartials_sum_571 ^ partials_44_14 ^
    partials_44_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_777 = reducedPartials_reducedPartials_sum_571 & partials_44_14 |
    partials_44_14 & partials_44_15 | reducedPartials_reducedPartials_sum_571 & partials_44_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_572 = reducedPartials_reducedPartials_carry_777 ^
    reducedPartials_reducedPartials_carry_776 ^ reducedPartials_reducedPartials_45_0_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_778 = reducedPartials_reducedPartials_carry_777 &
    reducedPartials_reducedPartials_carry_776 | reducedPartials_reducedPartials_carry_776 &
    reducedPartials_reducedPartials_45_0_3 | reducedPartials_reducedPartials_carry_777 &
    reducedPartials_reducedPartials_45_0_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_45_0_4 = reducedPartials_reducedPartials_sum_572 ^ partials_45_13 ^
    partials_45_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_779 = reducedPartials_reducedPartials_sum_572 & partials_45_13 |
    partials_45_13 & partials_45_14 | reducedPartials_reducedPartials_sum_572 & partials_45_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_573 = reducedPartials_reducedPartials_carry_779 ^
    reducedPartials_reducedPartials_carry_778 ^ reducedPartials_reducedPartials_46_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_780 = reducedPartials_reducedPartials_carry_779 &
    reducedPartials_reducedPartials_carry_778 | reducedPartials_reducedPartials_carry_778 &
    reducedPartials_reducedPartials_46_0_2 | reducedPartials_reducedPartials_carry_779 &
    reducedPartials_reducedPartials_46_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_46_0_3 = reducedPartials_reducedPartials_sum_573 ^ partials_46_12 ^
    partials_46_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_781 = reducedPartials_reducedPartials_sum_573 & partials_46_12 |
    partials_46_12 & partials_46_13 | reducedPartials_reducedPartials_sum_573 & partials_46_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_574 = reducedPartials_reducedPartials_carry_781 ^
    reducedPartials_reducedPartials_carry_780 ^ reducedPartials_reducedPartials_47_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_782 = reducedPartials_reducedPartials_carry_781 &
    reducedPartials_reducedPartials_carry_780 | reducedPartials_reducedPartials_carry_780 &
    reducedPartials_reducedPartials_47_0_2 | reducedPartials_reducedPartials_carry_781 &
    reducedPartials_reducedPartials_47_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_47_0_3 = reducedPartials_reducedPartials_sum_574 ^ partials_47_11 ^
    partials_47_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_783 = reducedPartials_reducedPartials_sum_574 & partials_47_11 |
    partials_47_11 & partials_47_12 | reducedPartials_reducedPartials_sum_574 & partials_47_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_575 = reducedPartials_reducedPartials_carry_783 ^
    reducedPartials_reducedPartials_carry_782 ^ reducedPartials_reducedPartials_48_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_784 = reducedPartials_reducedPartials_carry_783 &
    reducedPartials_reducedPartials_carry_782 | reducedPartials_reducedPartials_carry_782 &
    reducedPartials_reducedPartials_48_0_2 | reducedPartials_reducedPartials_carry_783 &
    reducedPartials_reducedPartials_48_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_48_0_3 = reducedPartials_reducedPartials_sum_575 ^ partials_48_10 ^
    partials_48_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_785 = reducedPartials_reducedPartials_sum_575 & partials_48_10 |
    partials_48_10 & partials_48_11 | reducedPartials_reducedPartials_sum_575 & partials_48_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_576 = reducedPartials_reducedPartials_carry_785 ^
    reducedPartials_reducedPartials_carry_784 ^ reducedPartials_reducedPartials_49_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_786 = reducedPartials_reducedPartials_carry_785 &
    reducedPartials_reducedPartials_carry_784 | reducedPartials_reducedPartials_carry_784 &
    reducedPartials_reducedPartials_49_0_2 | reducedPartials_reducedPartials_carry_785 &
    reducedPartials_reducedPartials_49_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_49_0_3 = reducedPartials_reducedPartials_sum_576 ^ partials_49_9 ^
    partials_49_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_787 = reducedPartials_reducedPartials_sum_576 & partials_49_9 |
    partials_49_9 & partials_49_10 | reducedPartials_reducedPartials_sum_576 & partials_49_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_577 = reducedPartials_reducedPartials_carry_787 ^
    reducedPartials_reducedPartials_carry_786 ^ reducedPartials_reducedPartials_50_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_788 = reducedPartials_reducedPartials_carry_787 &
    reducedPartials_reducedPartials_carry_786 | reducedPartials_reducedPartials_carry_786 &
    reducedPartials_reducedPartials_50_0_2 | reducedPartials_reducedPartials_carry_787 &
    reducedPartials_reducedPartials_50_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_50_0_3 = reducedPartials_reducedPartials_sum_577 ^ partials_50_8 ^ partials_50_9
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_789 = reducedPartials_reducedPartials_sum_577 & partials_50_8 |
    partials_50_8 & partials_50_9 | reducedPartials_reducedPartials_sum_577 & partials_50_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_578 = reducedPartials_reducedPartials_carry_789 ^
    reducedPartials_reducedPartials_carry_788 ^ reducedPartials_reducedPartials_51_0_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_790 = reducedPartials_reducedPartials_carry_789 &
    reducedPartials_reducedPartials_carry_788 | reducedPartials_reducedPartials_carry_788 &
    reducedPartials_reducedPartials_51_0_2 | reducedPartials_reducedPartials_carry_789 &
    reducedPartials_reducedPartials_51_0_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_51_0_3 = reducedPartials_reducedPartials_sum_578 ^ partials_51_7 ^ partials_51_8
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_791 = reducedPartials_reducedPartials_sum_578 & partials_51_7 |
    partials_51_7 & partials_51_8 | reducedPartials_reducedPartials_sum_578 & partials_51_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_579 = reducedPartials_reducedPartials_carry_791 ^
    reducedPartials_reducedPartials_carry_790 ^ reducedPartials_reducedPartials_52_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_792 = reducedPartials_reducedPartials_carry_791 &
    reducedPartials_reducedPartials_carry_790 | reducedPartials_reducedPartials_carry_790 &
    reducedPartials_reducedPartials_52_0_1 | reducedPartials_reducedPartials_carry_791 &
    reducedPartials_reducedPartials_52_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_52_0_2 = reducedPartials_reducedPartials_sum_579 ^ partials_52_6 ^ partials_52_7
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_793 = reducedPartials_reducedPartials_sum_579 & partials_52_6 |
    partials_52_6 & partials_52_7 | reducedPartials_reducedPartials_sum_579 & partials_52_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_580 = reducedPartials_reducedPartials_carry_793 ^
    reducedPartials_reducedPartials_carry_792 ^ reducedPartials_reducedPartials_53_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_794 = reducedPartials_reducedPartials_carry_793 &
    reducedPartials_reducedPartials_carry_792 | reducedPartials_reducedPartials_carry_792 &
    reducedPartials_reducedPartials_53_0_1 | reducedPartials_reducedPartials_carry_793 &
    reducedPartials_reducedPartials_53_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_53_0_2 = reducedPartials_reducedPartials_sum_580 ^ partials_53_5 ^ partials_53_6
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_795 = reducedPartials_reducedPartials_sum_580 & partials_53_5 |
    partials_53_5 & partials_53_6 | reducedPartials_reducedPartials_sum_580 & partials_53_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_581 = reducedPartials_reducedPartials_carry_795 ^
    reducedPartials_reducedPartials_carry_794 ^ reducedPartials_reducedPartials_54_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_796 = reducedPartials_reducedPartials_carry_795 &
    reducedPartials_reducedPartials_carry_794 | reducedPartials_reducedPartials_carry_794 &
    reducedPartials_reducedPartials_54_0_1 | reducedPartials_reducedPartials_carry_795 &
    reducedPartials_reducedPartials_54_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_54_0_2 = reducedPartials_reducedPartials_sum_581 ^ partials_54_4 ^ partials_54_5
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_797 = reducedPartials_reducedPartials_sum_581 & partials_54_4 |
    partials_54_4 & partials_54_5 | reducedPartials_reducedPartials_sum_581 & partials_54_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_582 = reducedPartials_reducedPartials_carry_797 ^
    reducedPartials_reducedPartials_carry_796 ^ reducedPartials_reducedPartials_55_0_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_798 = reducedPartials_reducedPartials_carry_797 &
    reducedPartials_reducedPartials_carry_796 | reducedPartials_reducedPartials_carry_796 &
    reducedPartials_reducedPartials_55_0_1 | reducedPartials_reducedPartials_carry_797 &
    reducedPartials_reducedPartials_55_0_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_55_0_2 = reducedPartials_reducedPartials_sum_582 ^ partials_55_3 ^ partials_55_4
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_799 = reducedPartials_reducedPartials_sum_582 & partials_55_3 |
    partials_55_3 & partials_55_4 | reducedPartials_reducedPartials_sum_582 & partials_55_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_583 = reducedPartials_reducedPartials_carry_799 ^
    reducedPartials_reducedPartials_carry_798 ^ reducedPartials_reducedPartials_56_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_800 = reducedPartials_reducedPartials_carry_799 &
    reducedPartials_reducedPartials_carry_798 | reducedPartials_reducedPartials_carry_798 &
    reducedPartials_reducedPartials_56_0 | reducedPartials_reducedPartials_carry_799 &
    reducedPartials_reducedPartials_56_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_56_0_1 = reducedPartials_reducedPartials_sum_583 ^ partials_56_2 ^ partials_56_3
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_801 = reducedPartials_reducedPartials_sum_583 & partials_56_2 |
    partials_56_2 & partials_56_3 | reducedPartials_reducedPartials_sum_583 & partials_56_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_584 = reducedPartials_reducedPartials_carry_801 ^
    reducedPartials_reducedPartials_carry_800 ^ reducedPartials_reducedPartials_57_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_802 = reducedPartials_reducedPartials_carry_801 &
    reducedPartials_reducedPartials_carry_800 | reducedPartials_reducedPartials_carry_800 &
    reducedPartials_reducedPartials_57_0 | reducedPartials_reducedPartials_carry_801 &
    reducedPartials_reducedPartials_57_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_57_0_1 = reducedPartials_reducedPartials_sum_584 ^ partials_57_1 ^ partials_57_2
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_803 = reducedPartials_reducedPartials_sum_584 & partials_57_1 |
    partials_57_1 & partials_57_2 | reducedPartials_reducedPartials_sum_584 & partials_57_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_sum_585 = reducedPartials_reducedPartials_carry_803 ^
    reducedPartials_reducedPartials_carry_802 ^ reducedPartials_reducedPartials_58_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_804 = reducedPartials_reducedPartials_carry_803 &
    reducedPartials_reducedPartials_carry_802 | reducedPartials_reducedPartials_carry_802 &
    reducedPartials_reducedPartials_58_0 | reducedPartials_reducedPartials_carry_803 &
    reducedPartials_reducedPartials_58_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_58_0_1 = reducedPartials_reducedPartials_sum_585 ^ partials_58_0 ^ partials_58_1
    ; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_805 = reducedPartials_reducedPartials_sum_585 & partials_58_0 |
    partials_58_0 & partials_58_1 | reducedPartials_reducedPartials_sum_585 & partials_58_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_59_0 = reducedPartials_reducedPartials_carry_805 ^
    reducedPartials_reducedPartials_carry_804 ^ partials_59_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_60_0 = reducedPartials_reducedPartials_carry_805 &
    reducedPartials_reducedPartials_carry_804 | reducedPartials_reducedPartials_carry_804 & partials_59_0 |
    reducedPartials_reducedPartials_carry_805 & partials_59_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_3_0 = partials_3_0 ^ partials_3_1; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_806 = partials_3_0 & partials_3_1; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_reducedPartials_4_0_1 = reducedPartials_reducedPartials_carry_806 ^
    reducedPartials_reducedPartials_4_0 ^ partials_4_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_807 = reducedPartials_reducedPartials_carry_806 &
    reducedPartials_reducedPartials_4_0 | reducedPartials_reducedPartials_4_0 & partials_4_2 |
    reducedPartials_reducedPartials_carry_806 & partials_4_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_5_0_1 = reducedPartials_reducedPartials_carry_807 ^
    reducedPartials_reducedPartials_5_0 ^ partials_5_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_808 = reducedPartials_reducedPartials_carry_807 &
    reducedPartials_reducedPartials_5_0 | reducedPartials_reducedPartials_5_0 & partials_5_3 |
    reducedPartials_reducedPartials_carry_807 & partials_5_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_6_0_2 = reducedPartials_reducedPartials_carry_808 ^
    reducedPartials_reducedPartials_6_0_1 ^ partials_6_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_809 = reducedPartials_reducedPartials_carry_808 &
    reducedPartials_reducedPartials_6_0_1 | reducedPartials_reducedPartials_6_0_1 & partials_6_4 |
    reducedPartials_reducedPartials_carry_808 & partials_6_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_7_0_2 = reducedPartials_reducedPartials_carry_809 ^
    reducedPartials_reducedPartials_7_0_1 ^ partials_7_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_810 = reducedPartials_reducedPartials_carry_809 &
    reducedPartials_reducedPartials_7_0_1 | reducedPartials_reducedPartials_7_0_1 & partials_7_5 |
    reducedPartials_reducedPartials_carry_809 & partials_7_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_8_0_2 = reducedPartials_reducedPartials_carry_810 ^
    reducedPartials_reducedPartials_8_0_1 ^ partials_8_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_811 = reducedPartials_reducedPartials_carry_810 &
    reducedPartials_reducedPartials_8_0_1 | reducedPartials_reducedPartials_8_0_1 & partials_8_6 |
    reducedPartials_reducedPartials_carry_810 & partials_8_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_9_0_3 = reducedPartials_reducedPartials_carry_811 ^
    reducedPartials_reducedPartials_9_0_2 ^ partials_9_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_812 = reducedPartials_reducedPartials_carry_811 &
    reducedPartials_reducedPartials_9_0_2 | reducedPartials_reducedPartials_9_0_2 & partials_9_7 |
    reducedPartials_reducedPartials_carry_811 & partials_9_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_10_0_3 = reducedPartials_reducedPartials_carry_812 ^
    reducedPartials_reducedPartials_10_0_2 ^ partials_10_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_813 = reducedPartials_reducedPartials_carry_812 &
    reducedPartials_reducedPartials_10_0_2 | reducedPartials_reducedPartials_10_0_2 & partials_10_8 |
    reducedPartials_reducedPartials_carry_812 & partials_10_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_11_0_3 = reducedPartials_reducedPartials_carry_813 ^
    reducedPartials_reducedPartials_11_0_2 ^ partials_11_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_814 = reducedPartials_reducedPartials_carry_813 &
    reducedPartials_reducedPartials_11_0_2 | reducedPartials_reducedPartials_11_0_2 & partials_11_9 |
    reducedPartials_reducedPartials_carry_813 & partials_11_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_12_0_3 = reducedPartials_reducedPartials_carry_814 ^
    reducedPartials_reducedPartials_12_0_2 ^ partials_12_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_815 = reducedPartials_reducedPartials_carry_814 &
    reducedPartials_reducedPartials_12_0_2 | reducedPartials_reducedPartials_12_0_2 & partials_12_10 |
    reducedPartials_reducedPartials_carry_814 & partials_12_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_13_0_4 = reducedPartials_reducedPartials_carry_815 ^
    reducedPartials_reducedPartials_13_0_3 ^ partials_13_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_816 = reducedPartials_reducedPartials_carry_815 &
    reducedPartials_reducedPartials_13_0_3 | reducedPartials_reducedPartials_13_0_3 & partials_13_11 |
    reducedPartials_reducedPartials_carry_815 & partials_13_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_14_0_4 = reducedPartials_reducedPartials_carry_816 ^
    reducedPartials_reducedPartials_14_0_3 ^ partials_14_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_817 = reducedPartials_reducedPartials_carry_816 &
    reducedPartials_reducedPartials_14_0_3 | reducedPartials_reducedPartials_14_0_3 & partials_14_12 |
    reducedPartials_reducedPartials_carry_816 & partials_14_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_15_0_4 = reducedPartials_reducedPartials_carry_817 ^
    reducedPartials_reducedPartials_15_0_3 ^ partials_15_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_818 = reducedPartials_reducedPartials_carry_817 &
    reducedPartials_reducedPartials_15_0_3 | reducedPartials_reducedPartials_15_0_3 & partials_15_13 |
    reducedPartials_reducedPartials_carry_817 & partials_15_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_16_0_4 = reducedPartials_reducedPartials_carry_818 ^
    reducedPartials_reducedPartials_16_0_3 ^ partials_16_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_819 = reducedPartials_reducedPartials_carry_818 &
    reducedPartials_reducedPartials_16_0_3 | reducedPartials_reducedPartials_16_0_3 & partials_16_14 |
    reducedPartials_reducedPartials_carry_818 & partials_16_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_17_0_4 = reducedPartials_reducedPartials_carry_819 ^
    reducedPartials_reducedPartials_17_0_3 ^ partials_17_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_820 = reducedPartials_reducedPartials_carry_819 &
    reducedPartials_reducedPartials_17_0_3 | reducedPartials_reducedPartials_17_0_3 & partials_17_15 |
    reducedPartials_reducedPartials_carry_819 & partials_17_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_18_0_4 = reducedPartials_reducedPartials_carry_820 ^
    reducedPartials_reducedPartials_18_0_3 ^ partials_18_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_821 = reducedPartials_reducedPartials_carry_820 &
    reducedPartials_reducedPartials_18_0_3 | reducedPartials_reducedPartials_18_0_3 & partials_18_16 |
    reducedPartials_reducedPartials_carry_820 & partials_18_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_19_0_5 = reducedPartials_reducedPartials_carry_821 ^
    reducedPartials_reducedPartials_19_0_4 ^ partials_19_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_822 = reducedPartials_reducedPartials_carry_821 &
    reducedPartials_reducedPartials_19_0_4 | reducedPartials_reducedPartials_19_0_4 & partials_19_17 |
    reducedPartials_reducedPartials_carry_821 & partials_19_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_20_0_5 = reducedPartials_reducedPartials_carry_822 ^
    reducedPartials_reducedPartials_20_0_4 ^ partials_20_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_823 = reducedPartials_reducedPartials_carry_822 &
    reducedPartials_reducedPartials_20_0_4 | reducedPartials_reducedPartials_20_0_4 & partials_20_18 |
    reducedPartials_reducedPartials_carry_822 & partials_20_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_21_0_5 = reducedPartials_reducedPartials_carry_823 ^
    reducedPartials_reducedPartials_21_0_4 ^ partials_21_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_824 = reducedPartials_reducedPartials_carry_823 &
    reducedPartials_reducedPartials_21_0_4 | reducedPartials_reducedPartials_21_0_4 & partials_21_19 |
    reducedPartials_reducedPartials_carry_823 & partials_21_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_22_0_5 = reducedPartials_reducedPartials_carry_824 ^
    reducedPartials_reducedPartials_22_0_4 ^ partials_22_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_825 = reducedPartials_reducedPartials_carry_824 &
    reducedPartials_reducedPartials_22_0_4 | reducedPartials_reducedPartials_22_0_4 & partials_22_20 |
    reducedPartials_reducedPartials_carry_824 & partials_22_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_23_0_5 = reducedPartials_reducedPartials_carry_825 ^
    reducedPartials_reducedPartials_23_0_4 ^ partials_23_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_826 = reducedPartials_reducedPartials_carry_825 &
    reducedPartials_reducedPartials_23_0_4 | reducedPartials_reducedPartials_23_0_4 & partials_23_21 |
    reducedPartials_reducedPartials_carry_825 & partials_23_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_24_0_5 = reducedPartials_reducedPartials_carry_826 ^
    reducedPartials_reducedPartials_24_0_4 ^ partials_24_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_827 = reducedPartials_reducedPartials_carry_826 &
    reducedPartials_reducedPartials_24_0_4 | reducedPartials_reducedPartials_24_0_4 & partials_24_22 |
    reducedPartials_reducedPartials_carry_826 & partials_24_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_25_0_5 = reducedPartials_reducedPartials_carry_827 ^
    reducedPartials_reducedPartials_25_0_4 ^ partials_25_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_828 = reducedPartials_reducedPartials_carry_827 &
    reducedPartials_reducedPartials_25_0_4 | reducedPartials_reducedPartials_25_0_4 & partials_25_23 |
    reducedPartials_reducedPartials_carry_827 & partials_25_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_26_0_5 = reducedPartials_reducedPartials_carry_828 ^
    reducedPartials_reducedPartials_26_0_4 ^ partials_26_24; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_829 = reducedPartials_reducedPartials_carry_828 &
    reducedPartials_reducedPartials_26_0_4 | reducedPartials_reducedPartials_26_0_4 & partials_26_24 |
    reducedPartials_reducedPartials_carry_828 & partials_26_24; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_27_0_5 = reducedPartials_reducedPartials_carry_829 ^
    reducedPartials_reducedPartials_27_0_4 ^ partials_27_25; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_830 = reducedPartials_reducedPartials_carry_829 &
    reducedPartials_reducedPartials_27_0_4 | reducedPartials_reducedPartials_27_0_4 & partials_27_25 |
    reducedPartials_reducedPartials_carry_829 & partials_27_25; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_28_0_6 = reducedPartials_reducedPartials_carry_830 ^
    reducedPartials_reducedPartials_28_0_5 ^ partials_28_26; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_831 = reducedPartials_reducedPartials_carry_830 &
    reducedPartials_reducedPartials_28_0_5 | reducedPartials_reducedPartials_28_0_5 & partials_28_26 |
    reducedPartials_reducedPartials_carry_830 & partials_28_26; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_29_0_6 = reducedPartials_reducedPartials_carry_831 ^
    reducedPartials_reducedPartials_29_0_5 ^ partials_29_27; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_832 = reducedPartials_reducedPartials_carry_831 &
    reducedPartials_reducedPartials_29_0_5 | reducedPartials_reducedPartials_29_0_5 & partials_29_27 |
    reducedPartials_reducedPartials_carry_831 & partials_29_27; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_30_0_6 = reducedPartials_reducedPartials_carry_832 ^
    reducedPartials_reducedPartials_30_0_5 ^ partials_30_28; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_833 = reducedPartials_reducedPartials_carry_832 &
    reducedPartials_reducedPartials_30_0_5 | reducedPartials_reducedPartials_30_0_5 & partials_30_28 |
    reducedPartials_reducedPartials_carry_832 & partials_30_28; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_31_0_6 = reducedPartials_reducedPartials_carry_833 ^
    reducedPartials_reducedPartials_31_0_5 ^ partials_31_29; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_834 = reducedPartials_reducedPartials_carry_833 &
    reducedPartials_reducedPartials_31_0_5 | reducedPartials_reducedPartials_31_0_5 & partials_31_29 |
    reducedPartials_reducedPartials_carry_833 & partials_31_29; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_32_0_6 = reducedPartials_reducedPartials_carry_834 ^
    reducedPartials_reducedPartials_32_0_5 ^ partials_32_28; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_835 = reducedPartials_reducedPartials_carry_834 &
    reducedPartials_reducedPartials_32_0_5 | reducedPartials_reducedPartials_32_0_5 & partials_32_28 |
    reducedPartials_reducedPartials_carry_834 & partials_32_28; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_33_0_6 = reducedPartials_reducedPartials_carry_835 ^
    reducedPartials_reducedPartials_33_0_5 ^ partials_33_27; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_836 = reducedPartials_reducedPartials_carry_835 &
    reducedPartials_reducedPartials_33_0_5 | reducedPartials_reducedPartials_33_0_5 & partials_33_27 |
    reducedPartials_reducedPartials_carry_835 & partials_33_27; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_34_0_6 = reducedPartials_reducedPartials_carry_836 ^
    reducedPartials_reducedPartials_34_0_5 ^ partials_34_26; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_837 = reducedPartials_reducedPartials_carry_836 &
    reducedPartials_reducedPartials_34_0_5 | reducedPartials_reducedPartials_34_0_5 & partials_34_26 |
    reducedPartials_reducedPartials_carry_836 & partials_34_26; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_35_0_6 = reducedPartials_reducedPartials_carry_837 ^
    reducedPartials_reducedPartials_35_0_5 ^ partials_35_25; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_838 = reducedPartials_reducedPartials_carry_837 &
    reducedPartials_reducedPartials_35_0_5 | reducedPartials_reducedPartials_35_0_5 & partials_35_25 |
    reducedPartials_reducedPartials_carry_837 & partials_35_25; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_36_0_6 = reducedPartials_reducedPartials_carry_838 ^
    reducedPartials_reducedPartials_36_0_5 ^ partials_36_24; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_839 = reducedPartials_reducedPartials_carry_838 &
    reducedPartials_reducedPartials_36_0_5 | reducedPartials_reducedPartials_36_0_5 & partials_36_24 |
    reducedPartials_reducedPartials_carry_838 & partials_36_24; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_37_0_5 = reducedPartials_reducedPartials_carry_839 ^
    reducedPartials_reducedPartials_37_0_4 ^ partials_37_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_840 = reducedPartials_reducedPartials_carry_839 &
    reducedPartials_reducedPartials_37_0_4 | reducedPartials_reducedPartials_37_0_4 & partials_37_23 |
    reducedPartials_reducedPartials_carry_839 & partials_37_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_38_0_5 = reducedPartials_reducedPartials_carry_840 ^
    reducedPartials_reducedPartials_38_0_4 ^ partials_38_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_841 = reducedPartials_reducedPartials_carry_840 &
    reducedPartials_reducedPartials_38_0_4 | reducedPartials_reducedPartials_38_0_4 & partials_38_22 |
    reducedPartials_reducedPartials_carry_840 & partials_38_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_39_0_5 = reducedPartials_reducedPartials_carry_841 ^
    reducedPartials_reducedPartials_39_0_4 ^ partials_39_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_842 = reducedPartials_reducedPartials_carry_841 &
    reducedPartials_reducedPartials_39_0_4 | reducedPartials_reducedPartials_39_0_4 & partials_39_21 |
    reducedPartials_reducedPartials_carry_841 & partials_39_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_40_0_5 = reducedPartials_reducedPartials_carry_842 ^
    reducedPartials_reducedPartials_40_0_4 ^ partials_40_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_843 = reducedPartials_reducedPartials_carry_842 &
    reducedPartials_reducedPartials_40_0_4 | reducedPartials_reducedPartials_40_0_4 & partials_40_20 |
    reducedPartials_reducedPartials_carry_842 & partials_40_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_41_0_5 = reducedPartials_reducedPartials_carry_843 ^
    reducedPartials_reducedPartials_41_0_4 ^ partials_41_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_844 = reducedPartials_reducedPartials_carry_843 &
    reducedPartials_reducedPartials_41_0_4 | reducedPartials_reducedPartials_41_0_4 & partials_41_19 |
    reducedPartials_reducedPartials_carry_843 & partials_41_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_42_0_5 = reducedPartials_reducedPartials_carry_844 ^
    reducedPartials_reducedPartials_42_0_4 ^ partials_42_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_845 = reducedPartials_reducedPartials_carry_844 &
    reducedPartials_reducedPartials_42_0_4 | reducedPartials_reducedPartials_42_0_4 & partials_42_18 |
    reducedPartials_reducedPartials_carry_844 & partials_42_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_43_0_5 = reducedPartials_reducedPartials_carry_845 ^
    reducedPartials_reducedPartials_43_0_4 ^ partials_43_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_846 = reducedPartials_reducedPartials_carry_845 &
    reducedPartials_reducedPartials_43_0_4 | reducedPartials_reducedPartials_43_0_4 & partials_43_17 |
    reducedPartials_reducedPartials_carry_845 & partials_43_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_44_0_5 = reducedPartials_reducedPartials_carry_846 ^
    reducedPartials_reducedPartials_44_0_4 ^ partials_44_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_847 = reducedPartials_reducedPartials_carry_846 &
    reducedPartials_reducedPartials_44_0_4 | reducedPartials_reducedPartials_44_0_4 & partials_44_16 |
    reducedPartials_reducedPartials_carry_846 & partials_44_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_45_0_5 = reducedPartials_reducedPartials_carry_847 ^
    reducedPartials_reducedPartials_45_0_4 ^ partials_45_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_848 = reducedPartials_reducedPartials_carry_847 &
    reducedPartials_reducedPartials_45_0_4 | reducedPartials_reducedPartials_45_0_4 & partials_45_15 |
    reducedPartials_reducedPartials_carry_847 & partials_45_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_46_0_4 = reducedPartials_reducedPartials_carry_848 ^
    reducedPartials_reducedPartials_46_0_3 ^ partials_46_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_849 = reducedPartials_reducedPartials_carry_848 &
    reducedPartials_reducedPartials_46_0_3 | reducedPartials_reducedPartials_46_0_3 & partials_46_14 |
    reducedPartials_reducedPartials_carry_848 & partials_46_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_47_0_4 = reducedPartials_reducedPartials_carry_849 ^
    reducedPartials_reducedPartials_47_0_3 ^ partials_47_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_850 = reducedPartials_reducedPartials_carry_849 &
    reducedPartials_reducedPartials_47_0_3 | reducedPartials_reducedPartials_47_0_3 & partials_47_13 |
    reducedPartials_reducedPartials_carry_849 & partials_47_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_48_0_4 = reducedPartials_reducedPartials_carry_850 ^
    reducedPartials_reducedPartials_48_0_3 ^ partials_48_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_851 = reducedPartials_reducedPartials_carry_850 &
    reducedPartials_reducedPartials_48_0_3 | reducedPartials_reducedPartials_48_0_3 & partials_48_12 |
    reducedPartials_reducedPartials_carry_850 & partials_48_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_49_0_4 = reducedPartials_reducedPartials_carry_851 ^
    reducedPartials_reducedPartials_49_0_3 ^ partials_49_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_852 = reducedPartials_reducedPartials_carry_851 &
    reducedPartials_reducedPartials_49_0_3 | reducedPartials_reducedPartials_49_0_3 & partials_49_11 |
    reducedPartials_reducedPartials_carry_851 & partials_49_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_50_0_4 = reducedPartials_reducedPartials_carry_852 ^
    reducedPartials_reducedPartials_50_0_3 ^ partials_50_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_853 = reducedPartials_reducedPartials_carry_852 &
    reducedPartials_reducedPartials_50_0_3 | reducedPartials_reducedPartials_50_0_3 & partials_50_10 |
    reducedPartials_reducedPartials_carry_852 & partials_50_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_51_0_4 = reducedPartials_reducedPartials_carry_853 ^
    reducedPartials_reducedPartials_51_0_3 ^ partials_51_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_854 = reducedPartials_reducedPartials_carry_853 &
    reducedPartials_reducedPartials_51_0_3 | reducedPartials_reducedPartials_51_0_3 & partials_51_9 |
    reducedPartials_reducedPartials_carry_853 & partials_51_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_52_0_3 = reducedPartials_reducedPartials_carry_854 ^
    reducedPartials_reducedPartials_52_0_2 ^ partials_52_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_855 = reducedPartials_reducedPartials_carry_854 &
    reducedPartials_reducedPartials_52_0_2 | reducedPartials_reducedPartials_52_0_2 & partials_52_8 |
    reducedPartials_reducedPartials_carry_854 & partials_52_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_53_0_3 = reducedPartials_reducedPartials_carry_855 ^
    reducedPartials_reducedPartials_53_0_2 ^ partials_53_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_856 = reducedPartials_reducedPartials_carry_855 &
    reducedPartials_reducedPartials_53_0_2 | reducedPartials_reducedPartials_53_0_2 & partials_53_7 |
    reducedPartials_reducedPartials_carry_855 & partials_53_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_54_0_3 = reducedPartials_reducedPartials_carry_856 ^
    reducedPartials_reducedPartials_54_0_2 ^ partials_54_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_857 = reducedPartials_reducedPartials_carry_856 &
    reducedPartials_reducedPartials_54_0_2 | reducedPartials_reducedPartials_54_0_2 & partials_54_6 |
    reducedPartials_reducedPartials_carry_856 & partials_54_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_55_0_3 = reducedPartials_reducedPartials_carry_857 ^
    reducedPartials_reducedPartials_55_0_2 ^ partials_55_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_858 = reducedPartials_reducedPartials_carry_857 &
    reducedPartials_reducedPartials_55_0_2 | reducedPartials_reducedPartials_55_0_2 & partials_55_5 |
    reducedPartials_reducedPartials_carry_857 & partials_55_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_56_0_2 = reducedPartials_reducedPartials_carry_858 ^
    reducedPartials_reducedPartials_56_0_1 ^ partials_56_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_859 = reducedPartials_reducedPartials_carry_858 &
    reducedPartials_reducedPartials_56_0_1 | reducedPartials_reducedPartials_56_0_1 & partials_56_4 |
    reducedPartials_reducedPartials_carry_858 & partials_56_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_57_0_2 = reducedPartials_reducedPartials_carry_859 ^
    reducedPartials_reducedPartials_57_0_1 ^ partials_57_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_860 = reducedPartials_reducedPartials_carry_859 &
    reducedPartials_reducedPartials_57_0_1 | reducedPartials_reducedPartials_57_0_1 & partials_57_3 |
    reducedPartials_reducedPartials_carry_859 & partials_57_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_58_0_2 = reducedPartials_reducedPartials_carry_860 ^
    reducedPartials_reducedPartials_58_0_1 ^ partials_58_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_861 = reducedPartials_reducedPartials_carry_860 &
    reducedPartials_reducedPartials_58_0_1 | reducedPartials_reducedPartials_58_0_1 & partials_58_2 |
    reducedPartials_reducedPartials_carry_860 & partials_58_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_59_0_1 = reducedPartials_reducedPartials_carry_861 ^
    reducedPartials_reducedPartials_59_0 ^ partials_59_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_862 = reducedPartials_reducedPartials_carry_861 &
    reducedPartials_reducedPartials_59_0 | reducedPartials_reducedPartials_59_0 & partials_59_1 |
    reducedPartials_reducedPartials_carry_861 & partials_59_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_reducedPartials_60_0_1 = reducedPartials_reducedPartials_carry_862 ^
    reducedPartials_reducedPartials_60_0 ^ partials_60_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_61_0 = reducedPartials_reducedPartials_carry_862 &
    reducedPartials_reducedPartials_60_0 | reducedPartials_reducedPartials_60_0 & partials_60_0 |
    reducedPartials_reducedPartials_carry_862 & partials_60_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_2_0 = partials_2_0 ^ partials_2_1; // @[src/main/scala/dadda_tree_mult.scala 109:15]
  wire  reducedPartials_reducedPartials_carry_863 = partials_2_0 & partials_2_1; // @[src/main/scala/dadda_tree_mult.scala 110:17]
  wire  reducedPartials_3_0 = reducedPartials_reducedPartials_carry_863 ^ reducedPartials_reducedPartials_3_0 ^
    partials_3_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_864 = reducedPartials_reducedPartials_carry_863 &
    reducedPartials_reducedPartials_3_0 | reducedPartials_reducedPartials_3_0 & partials_3_2 |
    reducedPartials_reducedPartials_carry_863 & partials_3_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_4_0 = reducedPartials_reducedPartials_carry_864 ^ reducedPartials_reducedPartials_4_0_1 ^
    partials_4_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_865 = reducedPartials_reducedPartials_carry_864 &
    reducedPartials_reducedPartials_4_0_1 | reducedPartials_reducedPartials_4_0_1 & partials_4_3 |
    reducedPartials_reducedPartials_carry_864 & partials_4_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_5_0 = reducedPartials_reducedPartials_carry_865 ^ reducedPartials_reducedPartials_5_0_1 ^
    partials_5_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_866 = reducedPartials_reducedPartials_carry_865 &
    reducedPartials_reducedPartials_5_0_1 | reducedPartials_reducedPartials_5_0_1 & partials_5_4 |
    reducedPartials_reducedPartials_carry_865 & partials_5_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_6_0 = reducedPartials_reducedPartials_carry_866 ^ reducedPartials_reducedPartials_6_0_2 ^
    partials_6_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_867 = reducedPartials_reducedPartials_carry_866 &
    reducedPartials_reducedPartials_6_0_2 | reducedPartials_reducedPartials_6_0_2 & partials_6_5 |
    reducedPartials_reducedPartials_carry_866 & partials_6_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_7_0 = reducedPartials_reducedPartials_carry_867 ^ reducedPartials_reducedPartials_7_0_2 ^
    partials_7_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_868 = reducedPartials_reducedPartials_carry_867 &
    reducedPartials_reducedPartials_7_0_2 | reducedPartials_reducedPartials_7_0_2 & partials_7_6 |
    reducedPartials_reducedPartials_carry_867 & partials_7_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_8_0 = reducedPartials_reducedPartials_carry_868 ^ reducedPartials_reducedPartials_8_0_2 ^
    partials_8_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_869 = reducedPartials_reducedPartials_carry_868 &
    reducedPartials_reducedPartials_8_0_2 | reducedPartials_reducedPartials_8_0_2 & partials_8_7 |
    reducedPartials_reducedPartials_carry_868 & partials_8_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_9_0 = reducedPartials_reducedPartials_carry_869 ^ reducedPartials_reducedPartials_9_0_3 ^
    partials_9_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_870 = reducedPartials_reducedPartials_carry_869 &
    reducedPartials_reducedPartials_9_0_3 | reducedPartials_reducedPartials_9_0_3 & partials_9_8 |
    reducedPartials_reducedPartials_carry_869 & partials_9_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_10_0 = reducedPartials_reducedPartials_carry_870 ^ reducedPartials_reducedPartials_10_0_3 ^
    partials_10_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_871 = reducedPartials_reducedPartials_carry_870 &
    reducedPartials_reducedPartials_10_0_3 | reducedPartials_reducedPartials_10_0_3 & partials_10_9 |
    reducedPartials_reducedPartials_carry_870 & partials_10_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_11_0 = reducedPartials_reducedPartials_carry_871 ^ reducedPartials_reducedPartials_11_0_3 ^
    partials_11_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_872 = reducedPartials_reducedPartials_carry_871 &
    reducedPartials_reducedPartials_11_0_3 | reducedPartials_reducedPartials_11_0_3 & partials_11_10 |
    reducedPartials_reducedPartials_carry_871 & partials_11_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_12_0 = reducedPartials_reducedPartials_carry_872 ^ reducedPartials_reducedPartials_12_0_3 ^
    partials_12_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_873 = reducedPartials_reducedPartials_carry_872 &
    reducedPartials_reducedPartials_12_0_3 | reducedPartials_reducedPartials_12_0_3 & partials_12_11 |
    reducedPartials_reducedPartials_carry_872 & partials_12_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_13_0 = reducedPartials_reducedPartials_carry_873 ^ reducedPartials_reducedPartials_13_0_4 ^
    partials_13_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_874 = reducedPartials_reducedPartials_carry_873 &
    reducedPartials_reducedPartials_13_0_4 | reducedPartials_reducedPartials_13_0_4 & partials_13_12 |
    reducedPartials_reducedPartials_carry_873 & partials_13_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_14_0 = reducedPartials_reducedPartials_carry_874 ^ reducedPartials_reducedPartials_14_0_4 ^
    partials_14_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_875 = reducedPartials_reducedPartials_carry_874 &
    reducedPartials_reducedPartials_14_0_4 | reducedPartials_reducedPartials_14_0_4 & partials_14_13 |
    reducedPartials_reducedPartials_carry_874 & partials_14_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_15_0 = reducedPartials_reducedPartials_carry_875 ^ reducedPartials_reducedPartials_15_0_4 ^
    partials_15_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_876 = reducedPartials_reducedPartials_carry_875 &
    reducedPartials_reducedPartials_15_0_4 | reducedPartials_reducedPartials_15_0_4 & partials_15_14 |
    reducedPartials_reducedPartials_carry_875 & partials_15_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_16_0 = reducedPartials_reducedPartials_carry_876 ^ reducedPartials_reducedPartials_16_0_4 ^
    partials_16_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_877 = reducedPartials_reducedPartials_carry_876 &
    reducedPartials_reducedPartials_16_0_4 | reducedPartials_reducedPartials_16_0_4 & partials_16_15 |
    reducedPartials_reducedPartials_carry_876 & partials_16_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_17_0 = reducedPartials_reducedPartials_carry_877 ^ reducedPartials_reducedPartials_17_0_4 ^
    partials_17_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_878 = reducedPartials_reducedPartials_carry_877 &
    reducedPartials_reducedPartials_17_0_4 | reducedPartials_reducedPartials_17_0_4 & partials_17_16 |
    reducedPartials_reducedPartials_carry_877 & partials_17_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_18_0 = reducedPartials_reducedPartials_carry_878 ^ reducedPartials_reducedPartials_18_0_4 ^
    partials_18_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_879 = reducedPartials_reducedPartials_carry_878 &
    reducedPartials_reducedPartials_18_0_4 | reducedPartials_reducedPartials_18_0_4 & partials_18_17 |
    reducedPartials_reducedPartials_carry_878 & partials_18_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_19_0 = reducedPartials_reducedPartials_carry_879 ^ reducedPartials_reducedPartials_19_0_5 ^
    partials_19_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_880 = reducedPartials_reducedPartials_carry_879 &
    reducedPartials_reducedPartials_19_0_5 | reducedPartials_reducedPartials_19_0_5 & partials_19_18 |
    reducedPartials_reducedPartials_carry_879 & partials_19_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_20_0 = reducedPartials_reducedPartials_carry_880 ^ reducedPartials_reducedPartials_20_0_5 ^
    partials_20_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_881 = reducedPartials_reducedPartials_carry_880 &
    reducedPartials_reducedPartials_20_0_5 | reducedPartials_reducedPartials_20_0_5 & partials_20_19 |
    reducedPartials_reducedPartials_carry_880 & partials_20_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_21_0 = reducedPartials_reducedPartials_carry_881 ^ reducedPartials_reducedPartials_21_0_5 ^
    partials_21_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_882 = reducedPartials_reducedPartials_carry_881 &
    reducedPartials_reducedPartials_21_0_5 | reducedPartials_reducedPartials_21_0_5 & partials_21_20 |
    reducedPartials_reducedPartials_carry_881 & partials_21_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_22_0 = reducedPartials_reducedPartials_carry_882 ^ reducedPartials_reducedPartials_22_0_5 ^
    partials_22_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_883 = reducedPartials_reducedPartials_carry_882 &
    reducedPartials_reducedPartials_22_0_5 | reducedPartials_reducedPartials_22_0_5 & partials_22_21 |
    reducedPartials_reducedPartials_carry_882 & partials_22_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_23_0 = reducedPartials_reducedPartials_carry_883 ^ reducedPartials_reducedPartials_23_0_5 ^
    partials_23_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_884 = reducedPartials_reducedPartials_carry_883 &
    reducedPartials_reducedPartials_23_0_5 | reducedPartials_reducedPartials_23_0_5 & partials_23_22 |
    reducedPartials_reducedPartials_carry_883 & partials_23_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_24_0 = reducedPartials_reducedPartials_carry_884 ^ reducedPartials_reducedPartials_24_0_5 ^
    partials_24_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_885 = reducedPartials_reducedPartials_carry_884 &
    reducedPartials_reducedPartials_24_0_5 | reducedPartials_reducedPartials_24_0_5 & partials_24_23 |
    reducedPartials_reducedPartials_carry_884 & partials_24_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_25_0 = reducedPartials_reducedPartials_carry_885 ^ reducedPartials_reducedPartials_25_0_5 ^
    partials_25_24; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_886 = reducedPartials_reducedPartials_carry_885 &
    reducedPartials_reducedPartials_25_0_5 | reducedPartials_reducedPartials_25_0_5 & partials_25_24 |
    reducedPartials_reducedPartials_carry_885 & partials_25_24; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_26_0 = reducedPartials_reducedPartials_carry_886 ^ reducedPartials_reducedPartials_26_0_5 ^
    partials_26_25; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_887 = reducedPartials_reducedPartials_carry_886 &
    reducedPartials_reducedPartials_26_0_5 | reducedPartials_reducedPartials_26_0_5 & partials_26_25 |
    reducedPartials_reducedPartials_carry_886 & partials_26_25; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_27_0 = reducedPartials_reducedPartials_carry_887 ^ reducedPartials_reducedPartials_27_0_5 ^
    partials_27_26; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_888 = reducedPartials_reducedPartials_carry_887 &
    reducedPartials_reducedPartials_27_0_5 | reducedPartials_reducedPartials_27_0_5 & partials_27_26 |
    reducedPartials_reducedPartials_carry_887 & partials_27_26; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_28_0 = reducedPartials_reducedPartials_carry_888 ^ reducedPartials_reducedPartials_28_0_6 ^
    partials_28_27; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_889 = reducedPartials_reducedPartials_carry_888 &
    reducedPartials_reducedPartials_28_0_6 | reducedPartials_reducedPartials_28_0_6 & partials_28_27 |
    reducedPartials_reducedPartials_carry_888 & partials_28_27; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_29_0 = reducedPartials_reducedPartials_carry_889 ^ reducedPartials_reducedPartials_29_0_6 ^
    partials_29_28; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_890 = reducedPartials_reducedPartials_carry_889 &
    reducedPartials_reducedPartials_29_0_6 | reducedPartials_reducedPartials_29_0_6 & partials_29_28 |
    reducedPartials_reducedPartials_carry_889 & partials_29_28; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_30_0 = reducedPartials_reducedPartials_carry_890 ^ reducedPartials_reducedPartials_30_0_6 ^
    partials_30_29; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_891 = reducedPartials_reducedPartials_carry_890 &
    reducedPartials_reducedPartials_30_0_6 | reducedPartials_reducedPartials_30_0_6 & partials_30_29 |
    reducedPartials_reducedPartials_carry_890 & partials_30_29; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_31_0 = reducedPartials_reducedPartials_carry_891 ^ reducedPartials_reducedPartials_31_0_6 ^
    partials_31_30; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_892 = reducedPartials_reducedPartials_carry_891 &
    reducedPartials_reducedPartials_31_0_6 | reducedPartials_reducedPartials_31_0_6 & partials_31_30 |
    reducedPartials_reducedPartials_carry_891 & partials_31_30; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_32_0 = reducedPartials_reducedPartials_carry_892 ^ reducedPartials_reducedPartials_32_0_6 ^
    partials_32_29; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_893 = reducedPartials_reducedPartials_carry_892 &
    reducedPartials_reducedPartials_32_0_6 | reducedPartials_reducedPartials_32_0_6 & partials_32_29 |
    reducedPartials_reducedPartials_carry_892 & partials_32_29; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_33_0 = reducedPartials_reducedPartials_carry_893 ^ reducedPartials_reducedPartials_33_0_6 ^
    partials_33_28; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_894 = reducedPartials_reducedPartials_carry_893 &
    reducedPartials_reducedPartials_33_0_6 | reducedPartials_reducedPartials_33_0_6 & partials_33_28 |
    reducedPartials_reducedPartials_carry_893 & partials_33_28; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_34_0 = reducedPartials_reducedPartials_carry_894 ^ reducedPartials_reducedPartials_34_0_6 ^
    partials_34_27; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_895 = reducedPartials_reducedPartials_carry_894 &
    reducedPartials_reducedPartials_34_0_6 | reducedPartials_reducedPartials_34_0_6 & partials_34_27 |
    reducedPartials_reducedPartials_carry_894 & partials_34_27; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_35_0 = reducedPartials_reducedPartials_carry_895 ^ reducedPartials_reducedPartials_35_0_6 ^
    partials_35_26; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_896 = reducedPartials_reducedPartials_carry_895 &
    reducedPartials_reducedPartials_35_0_6 | reducedPartials_reducedPartials_35_0_6 & partials_35_26 |
    reducedPartials_reducedPartials_carry_895 & partials_35_26; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_36_0 = reducedPartials_reducedPartials_carry_896 ^ reducedPartials_reducedPartials_36_0_6 ^
    partials_36_25; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_897 = reducedPartials_reducedPartials_carry_896 &
    reducedPartials_reducedPartials_36_0_6 | reducedPartials_reducedPartials_36_0_6 & partials_36_25 |
    reducedPartials_reducedPartials_carry_896 & partials_36_25; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_37_0 = reducedPartials_reducedPartials_carry_897 ^ reducedPartials_reducedPartials_37_0_5 ^
    partials_37_24; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_898 = reducedPartials_reducedPartials_carry_897 &
    reducedPartials_reducedPartials_37_0_5 | reducedPartials_reducedPartials_37_0_5 & partials_37_24 |
    reducedPartials_reducedPartials_carry_897 & partials_37_24; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_38_0 = reducedPartials_reducedPartials_carry_898 ^ reducedPartials_reducedPartials_38_0_5 ^
    partials_38_23; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_899 = reducedPartials_reducedPartials_carry_898 &
    reducedPartials_reducedPartials_38_0_5 | reducedPartials_reducedPartials_38_0_5 & partials_38_23 |
    reducedPartials_reducedPartials_carry_898 & partials_38_23; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_39_0 = reducedPartials_reducedPartials_carry_899 ^ reducedPartials_reducedPartials_39_0_5 ^
    partials_39_22; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_900 = reducedPartials_reducedPartials_carry_899 &
    reducedPartials_reducedPartials_39_0_5 | reducedPartials_reducedPartials_39_0_5 & partials_39_22 |
    reducedPartials_reducedPartials_carry_899 & partials_39_22; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_40_0 = reducedPartials_reducedPartials_carry_900 ^ reducedPartials_reducedPartials_40_0_5 ^
    partials_40_21; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_901 = reducedPartials_reducedPartials_carry_900 &
    reducedPartials_reducedPartials_40_0_5 | reducedPartials_reducedPartials_40_0_5 & partials_40_21 |
    reducedPartials_reducedPartials_carry_900 & partials_40_21; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_41_0 = reducedPartials_reducedPartials_carry_901 ^ reducedPartials_reducedPartials_41_0_5 ^
    partials_41_20; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_902 = reducedPartials_reducedPartials_carry_901 &
    reducedPartials_reducedPartials_41_0_5 | reducedPartials_reducedPartials_41_0_5 & partials_41_20 |
    reducedPartials_reducedPartials_carry_901 & partials_41_20; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_42_0 = reducedPartials_reducedPartials_carry_902 ^ reducedPartials_reducedPartials_42_0_5 ^
    partials_42_19; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_903 = reducedPartials_reducedPartials_carry_902 &
    reducedPartials_reducedPartials_42_0_5 | reducedPartials_reducedPartials_42_0_5 & partials_42_19 |
    reducedPartials_reducedPartials_carry_902 & partials_42_19; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_43_0 = reducedPartials_reducedPartials_carry_903 ^ reducedPartials_reducedPartials_43_0_5 ^
    partials_43_18; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_904 = reducedPartials_reducedPartials_carry_903 &
    reducedPartials_reducedPartials_43_0_5 | reducedPartials_reducedPartials_43_0_5 & partials_43_18 |
    reducedPartials_reducedPartials_carry_903 & partials_43_18; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_44_0 = reducedPartials_reducedPartials_carry_904 ^ reducedPartials_reducedPartials_44_0_5 ^
    partials_44_17; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_905 = reducedPartials_reducedPartials_carry_904 &
    reducedPartials_reducedPartials_44_0_5 | reducedPartials_reducedPartials_44_0_5 & partials_44_17 |
    reducedPartials_reducedPartials_carry_904 & partials_44_17; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_45_0 = reducedPartials_reducedPartials_carry_905 ^ reducedPartials_reducedPartials_45_0_5 ^
    partials_45_16; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_906 = reducedPartials_reducedPartials_carry_905 &
    reducedPartials_reducedPartials_45_0_5 | reducedPartials_reducedPartials_45_0_5 & partials_45_16 |
    reducedPartials_reducedPartials_carry_905 & partials_45_16; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_46_0 = reducedPartials_reducedPartials_carry_906 ^ reducedPartials_reducedPartials_46_0_4 ^
    partials_46_15; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_907 = reducedPartials_reducedPartials_carry_906 &
    reducedPartials_reducedPartials_46_0_4 | reducedPartials_reducedPartials_46_0_4 & partials_46_15 |
    reducedPartials_reducedPartials_carry_906 & partials_46_15; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_47_0 = reducedPartials_reducedPartials_carry_907 ^ reducedPartials_reducedPartials_47_0_4 ^
    partials_47_14; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_908 = reducedPartials_reducedPartials_carry_907 &
    reducedPartials_reducedPartials_47_0_4 | reducedPartials_reducedPartials_47_0_4 & partials_47_14 |
    reducedPartials_reducedPartials_carry_907 & partials_47_14; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_48_0 = reducedPartials_reducedPartials_carry_908 ^ reducedPartials_reducedPartials_48_0_4 ^
    partials_48_13; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_909 = reducedPartials_reducedPartials_carry_908 &
    reducedPartials_reducedPartials_48_0_4 | reducedPartials_reducedPartials_48_0_4 & partials_48_13 |
    reducedPartials_reducedPartials_carry_908 & partials_48_13; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_49_0 = reducedPartials_reducedPartials_carry_909 ^ reducedPartials_reducedPartials_49_0_4 ^
    partials_49_12; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_910 = reducedPartials_reducedPartials_carry_909 &
    reducedPartials_reducedPartials_49_0_4 | reducedPartials_reducedPartials_49_0_4 & partials_49_12 |
    reducedPartials_reducedPartials_carry_909 & partials_49_12; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_50_0 = reducedPartials_reducedPartials_carry_910 ^ reducedPartials_reducedPartials_50_0_4 ^
    partials_50_11; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_911 = reducedPartials_reducedPartials_carry_910 &
    reducedPartials_reducedPartials_50_0_4 | reducedPartials_reducedPartials_50_0_4 & partials_50_11 |
    reducedPartials_reducedPartials_carry_910 & partials_50_11; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_51_0 = reducedPartials_reducedPartials_carry_911 ^ reducedPartials_reducedPartials_51_0_4 ^
    partials_51_10; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_912 = reducedPartials_reducedPartials_carry_911 &
    reducedPartials_reducedPartials_51_0_4 | reducedPartials_reducedPartials_51_0_4 & partials_51_10 |
    reducedPartials_reducedPartials_carry_911 & partials_51_10; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_52_0 = reducedPartials_reducedPartials_carry_912 ^ reducedPartials_reducedPartials_52_0_3 ^
    partials_52_9; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_913 = reducedPartials_reducedPartials_carry_912 &
    reducedPartials_reducedPartials_52_0_3 | reducedPartials_reducedPartials_52_0_3 & partials_52_9 |
    reducedPartials_reducedPartials_carry_912 & partials_52_9; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_53_0 = reducedPartials_reducedPartials_carry_913 ^ reducedPartials_reducedPartials_53_0_3 ^
    partials_53_8; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_914 = reducedPartials_reducedPartials_carry_913 &
    reducedPartials_reducedPartials_53_0_3 | reducedPartials_reducedPartials_53_0_3 & partials_53_8 |
    reducedPartials_reducedPartials_carry_913 & partials_53_8; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_54_0 = reducedPartials_reducedPartials_carry_914 ^ reducedPartials_reducedPartials_54_0_3 ^
    partials_54_7; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_915 = reducedPartials_reducedPartials_carry_914 &
    reducedPartials_reducedPartials_54_0_3 | reducedPartials_reducedPartials_54_0_3 & partials_54_7 |
    reducedPartials_reducedPartials_carry_914 & partials_54_7; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_55_0 = reducedPartials_reducedPartials_carry_915 ^ reducedPartials_reducedPartials_55_0_3 ^
    partials_55_6; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_916 = reducedPartials_reducedPartials_carry_915 &
    reducedPartials_reducedPartials_55_0_3 | reducedPartials_reducedPartials_55_0_3 & partials_55_6 |
    reducedPartials_reducedPartials_carry_915 & partials_55_6; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_56_0 = reducedPartials_reducedPartials_carry_916 ^ reducedPartials_reducedPartials_56_0_2 ^
    partials_56_5; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_917 = reducedPartials_reducedPartials_carry_916 &
    reducedPartials_reducedPartials_56_0_2 | reducedPartials_reducedPartials_56_0_2 & partials_56_5 |
    reducedPartials_reducedPartials_carry_916 & partials_56_5; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_57_0 = reducedPartials_reducedPartials_carry_917 ^ reducedPartials_reducedPartials_57_0_2 ^
    partials_57_4; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_918 = reducedPartials_reducedPartials_carry_917 &
    reducedPartials_reducedPartials_57_0_2 | reducedPartials_reducedPartials_57_0_2 & partials_57_4 |
    reducedPartials_reducedPartials_carry_917 & partials_57_4; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_58_0 = reducedPartials_reducedPartials_carry_918 ^ reducedPartials_reducedPartials_58_0_2 ^
    partials_58_3; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_919 = reducedPartials_reducedPartials_carry_918 &
    reducedPartials_reducedPartials_58_0_2 | reducedPartials_reducedPartials_58_0_2 & partials_58_3 |
    reducedPartials_reducedPartials_carry_918 & partials_58_3; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_59_0 = reducedPartials_reducedPartials_carry_919 ^ reducedPartials_reducedPartials_59_0_1 ^
    partials_59_2; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_920 = reducedPartials_reducedPartials_carry_919 &
    reducedPartials_reducedPartials_59_0_1 | reducedPartials_reducedPartials_59_0_1 & partials_59_2 |
    reducedPartials_reducedPartials_carry_919 & partials_59_2; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_60_0 = reducedPartials_reducedPartials_carry_920 ^ reducedPartials_reducedPartials_60_0_1 ^
    partials_60_1; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_reducedPartials_carry_921 = reducedPartials_reducedPartials_carry_920 &
    reducedPartials_reducedPartials_60_0_1 | reducedPartials_reducedPartials_60_0_1 & partials_60_1 |
    reducedPartials_reducedPartials_carry_920 & partials_60_1; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire  reducedPartials_61_0 = reducedPartials_reducedPartials_carry_921 ^ reducedPartials_reducedPartials_61_0 ^
    partials_61_0; // @[src/main/scala/dadda_tree_mult.scala 103:19]
  wire  reducedPartials_62_0 = reducedPartials_reducedPartials_carry_921 & reducedPartials_reducedPartials_61_0 |
    reducedPartials_reducedPartials_61_0 & partials_61_0 | reducedPartials_reducedPartials_carry_921 & partials_61_0; // @[src/main/scala/dadda_tree_mult.scala 104:35]
  wire [6:0] io_product_lo_lo_lo = {reducedPartials_6_0,reducedPartials_5_0,reducedPartials_4_0,reducedPartials_3_0,
    reducedPartials_2_0,partials_1_0,partials_0_0}; // @[src/main/scala/dadda_tree_mult.scala 162:28]
  wire [14:0] io_product_lo_lo = {reducedPartials_14_0,reducedPartials_13_0,reducedPartials_12_0,reducedPartials_11_0,
    reducedPartials_10_0,reducedPartials_9_0,reducedPartials_8_0,reducedPartials_7_0,io_product_lo_lo_lo}; // @[src/main/scala/dadda_tree_mult.scala 162:28]
  wire [7:0] io_product_lo_hi_lo = {reducedPartials_22_0,reducedPartials_21_0,reducedPartials_20_0,reducedPartials_19_0,
    reducedPartials_18_0,reducedPartials_17_0,reducedPartials_16_0,reducedPartials_15_0}; // @[src/main/scala/dadda_tree_mult.scala 162:28]
  wire [30:0] io_product_lo = {reducedPartials_30_0,reducedPartials_29_0,reducedPartials_28_0,reducedPartials_27_0,
    reducedPartials_26_0,reducedPartials_25_0,reducedPartials_24_0,reducedPartials_23_0,io_product_lo_hi_lo,
    io_product_lo_lo}; // @[src/main/scala/dadda_tree_mult.scala 162:28]
  wire [7:0] io_product_hi_lo_lo = {reducedPartials_38_0,reducedPartials_37_0,reducedPartials_36_0,reducedPartials_35_0,
    reducedPartials_34_0,reducedPartials_33_0,reducedPartials_32_0,reducedPartials_31_0}; // @[src/main/scala/dadda_tree_mult.scala 162:28]
  wire [15:0] io_product_hi_lo = {reducedPartials_46_0,reducedPartials_45_0,reducedPartials_44_0,reducedPartials_43_0,
    reducedPartials_42_0,reducedPartials_41_0,reducedPartials_40_0,reducedPartials_39_0,io_product_hi_lo_lo}; // @[src/main/scala/dadda_tree_mult.scala 162:28]
  wire [7:0] io_product_hi_hi_lo = {reducedPartials_54_0,reducedPartials_53_0,reducedPartials_52_0,reducedPartials_51_0,
    reducedPartials_50_0,reducedPartials_49_0,reducedPartials_48_0,reducedPartials_47_0}; // @[src/main/scala/dadda_tree_mult.scala 162:28]
  wire [31:0] io_product_hi = {reducedPartials_62_0,reducedPartials_61_0,reducedPartials_60_0,reducedPartials_59_0,
    reducedPartials_58_0,reducedPartials_57_0,reducedPartials_56_0,reducedPartials_55_0,io_product_hi_hi_lo,
    io_product_hi_lo}; // @[src/main/scala/dadda_tree_mult.scala 162:28]
  wire [6:0] io_product_lo_lo_lo_1 = {partials_6_6,partials_5_5,partials_4_4,partials_3_3,partials_2_2,partials_1_1,1'h0
    }; // @[src/main/scala/dadda_tree_mult.scala 162:48]
  wire [14:0] io_product_lo_lo_1 = {partials_14_14,partials_13_13,partials_12_12,partials_11_11,partials_10_10,
    partials_9_9,partials_8_8,partials_7_7,io_product_lo_lo_lo_1}; // @[src/main/scala/dadda_tree_mult.scala 162:48]
  wire [7:0] io_product_lo_hi_lo_1 = {partials_22_22,partials_21_21,partials_20_20,partials_19_19,partials_18_18,
    partials_17_17,partials_16_16,partials_15_15}; // @[src/main/scala/dadda_tree_mult.scala 162:48]
  wire [30:0] io_product_lo_1 = {partials_30_30,partials_29_29,partials_28_28,partials_27_27,partials_26_26,
    partials_25_25,partials_24_24,partials_23_23,io_product_lo_hi_lo_1,io_product_lo_lo_1}; // @[src/main/scala/dadda_tree_mult.scala 162:48]
  wire [7:0] io_product_hi_lo_lo_1 = {partials_38_24,partials_37_25,partials_36_26,partials_35_27,partials_34_28,
    partials_33_29,partials_32_30,partials_31_31}; // @[src/main/scala/dadda_tree_mult.scala 162:48]
  wire [15:0] io_product_hi_lo_1 = {partials_46_16,partials_45_17,partials_44_18,partials_43_19,partials_42_20,
    partials_41_21,partials_40_22,partials_39_23,io_product_hi_lo_lo_1}; // @[src/main/scala/dadda_tree_mult.scala 162:48]
  wire [7:0] io_product_hi_hi_lo_1 = {partials_54_8,partials_53_9,partials_52_10,partials_51_11,partials_50_12,
    partials_49_13,partials_48_14,partials_47_15}; // @[src/main/scala/dadda_tree_mult.scala 162:48]
  wire [31:0] io_product_hi_1 = {partials_62_0,partials_61_1,partials_60_2,partials_59_3,partials_58_4,partials_57_5,
    partials_56_6,partials_55_7,io_product_hi_hi_lo_1,io_product_hi_lo_1}; // @[src/main/scala/dadda_tree_mult.scala 162:48]
  RippleCarryAdder io_product_rca ( // @[src/main/scala/dadda_tree_mult.scala 163:21]
    .io_a(io_product_rca_io_a),
    .io_b(io_product_rca_io_b),
    .io_sum(io_product_rca_io_sum),
    .io_cout(io_product_rca_io_cout)
  );
  assign io_product = {io_product_rca_io_cout,io_product_rca_io_sum}; // @[src/main/scala/dadda_tree_mult.scala 168:8]
  assign io_product_rca_io_a = {io_product_hi,io_product_lo}; // @[src/main/scala/dadda_tree_mult.scala 162:28]
  assign io_product_rca_io_b = {io_product_hi_1,io_product_lo_1}; // @[src/main/scala/dadda_tree_mult.scala 162:48]
endmodule
