VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DaddaTreeMultiplier
  CLASS BLOCK ;
  FOREIGN DaddaTreeMultiplier ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 1756.000 700.030 1760.000 ;
    END
  END clock
  PIN io_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 35.400 2800.000 36.000 ;
    END
  END io_a[0]
  PIN io_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 579.400 2800.000 580.000 ;
    END
  END io_a[10]
  PIN io_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 633.800 2800.000 634.400 ;
    END
  END io_a[11]
  PIN io_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 688.200 2800.000 688.800 ;
    END
  END io_a[12]
  PIN io_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 742.600 2800.000 743.200 ;
    END
  END io_a[13]
  PIN io_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 797.000 2800.000 797.600 ;
    END
  END io_a[14]
  PIN io_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 851.400 2800.000 852.000 ;
    END
  END io_a[15]
  PIN io_a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 905.800 2800.000 906.400 ;
    END
  END io_a[16]
  PIN io_a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 960.200 2800.000 960.800 ;
    END
  END io_a[17]
  PIN io_a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1014.600 2800.000 1015.200 ;
    END
  END io_a[18]
  PIN io_a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1069.000 2800.000 1069.600 ;
    END
  END io_a[19]
  PIN io_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 89.800 2800.000 90.400 ;
    END
  END io_a[1]
  PIN io_a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1123.400 2800.000 1124.000 ;
    END
  END io_a[20]
  PIN io_a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1177.800 2800.000 1178.400 ;
    END
  END io_a[21]
  PIN io_a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1232.200 2800.000 1232.800 ;
    END
  END io_a[22]
  PIN io_a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1286.600 2800.000 1287.200 ;
    END
  END io_a[23]
  PIN io_a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1341.000 2800.000 1341.600 ;
    END
  END io_a[24]
  PIN io_a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1395.400 2800.000 1396.000 ;
    END
  END io_a[25]
  PIN io_a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1449.800 2800.000 1450.400 ;
    END
  END io_a[26]
  PIN io_a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1504.200 2800.000 1504.800 ;
    END
  END io_a[27]
  PIN io_a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1558.600 2800.000 1559.200 ;
    END
  END io_a[28]
  PIN io_a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1613.000 2800.000 1613.600 ;
    END
  END io_a[29]
  PIN io_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 144.200 2800.000 144.800 ;
    END
  END io_a[2]
  PIN io_a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1667.400 2800.000 1668.000 ;
    END
  END io_a[30]
  PIN io_a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1721.800 2800.000 1722.400 ;
    END
  END io_a[31]
  PIN io_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 198.600 2800.000 199.200 ;
    END
  END io_a[3]
  PIN io_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 253.000 2800.000 253.600 ;
    END
  END io_a[4]
  PIN io_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 307.400 2800.000 308.000 ;
    END
  END io_a[5]
  PIN io_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 361.800 2800.000 362.400 ;
    END
  END io_a[6]
  PIN io_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 416.200 2800.000 416.800 ;
    END
  END io_a[7]
  PIN io_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 470.600 2800.000 471.200 ;
    END
  END io_a[8]
  PIN io_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 525.000 2800.000 525.600 ;
    END
  END io_a[9]
  PIN io_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_b[0]
  PIN io_b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END io_b[10]
  PIN io_b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END io_b[11]
  PIN io_b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END io_b[12]
  PIN io_b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 742.600 4.000 743.200 ;
    END
  END io_b[13]
  PIN io_b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END io_b[14]
  PIN io_b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 4.000 852.000 ;
    END
  END io_b[15]
  PIN io_b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END io_b[16]
  PIN io_b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.200 4.000 960.800 ;
    END
  END io_b[17]
  PIN io_b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1014.600 4.000 1015.200 ;
    END
  END io_b[18]
  PIN io_b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1069.000 4.000 1069.600 ;
    END
  END io_b[19]
  PIN io_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_b[1]
  PIN io_b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1123.400 4.000 1124.000 ;
    END
  END io_b[20]
  PIN io_b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.800 4.000 1178.400 ;
    END
  END io_b[21]
  PIN io_b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1232.200 4.000 1232.800 ;
    END
  END io_b[22]
  PIN io_b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1286.600 4.000 1287.200 ;
    END
  END io_b[23]
  PIN io_b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1341.000 4.000 1341.600 ;
    END
  END io_b[24]
  PIN io_b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1395.400 4.000 1396.000 ;
    END
  END io_b[25]
  PIN io_b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1449.800 4.000 1450.400 ;
    END
  END io_b[26]
  PIN io_b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1504.200 4.000 1504.800 ;
    END
  END io_b[27]
  PIN io_b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1558.600 4.000 1559.200 ;
    END
  END io_b[28]
  PIN io_b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1613.000 4.000 1613.600 ;
    END
  END io_b[29]
  PIN io_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END io_b[2]
  PIN io_b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1667.400 4.000 1668.000 ;
    END
  END io_b[30]
  PIN io_b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1721.800 4.000 1722.400 ;
    END
  END io_b[31]
  PIN io_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END io_b[3]
  PIN io_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END io_b[4]
  PIN io_b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END io_b[5]
  PIN io_b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END io_b[6]
  PIN io_b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END io_b[7]
  PIN io_b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END io_b[8]
  PIN io_b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END io_b[9]
  PIN io_product[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END io_product[0]
  PIN io_product[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END io_product[10]
  PIN io_product[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END io_product[11]
  PIN io_product[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END io_product[12]
  PIN io_product[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END io_product[13]
  PIN io_product[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END io_product[14]
  PIN io_product[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END io_product[15]
  PIN io_product[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END io_product[16]
  PIN io_product[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END io_product[17]
  PIN io_product[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END io_product[18]
  PIN io_product[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END io_product[19]
  PIN io_product[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END io_product[1]
  PIN io_product[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 897.090 0.000 897.370 4.000 ;
    END
  END io_product[20]
  PIN io_product[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 940.790 0.000 941.070 4.000 ;
    END
  END io_product[21]
  PIN io_product[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 984.490 0.000 984.770 4.000 ;
    END
  END io_product[22]
  PIN io_product[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1028.190 0.000 1028.470 4.000 ;
    END
  END io_product[23]
  PIN io_product[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 4.000 ;
    END
  END io_product[24]
  PIN io_product[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1115.590 0.000 1115.870 4.000 ;
    END
  END io_product[25]
  PIN io_product[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END io_product[26]
  PIN io_product[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1202.990 0.000 1203.270 4.000 ;
    END
  END io_product[27]
  PIN io_product[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1246.690 0.000 1246.970 4.000 ;
    END
  END io_product[28]
  PIN io_product[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1290.390 0.000 1290.670 4.000 ;
    END
  END io_product[29]
  PIN io_product[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END io_product[2]
  PIN io_product[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1334.090 0.000 1334.370 4.000 ;
    END
  END io_product[30]
  PIN io_product[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1377.790 0.000 1378.070 4.000 ;
    END
  END io_product[31]
  PIN io_product[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1421.490 0.000 1421.770 4.000 ;
    END
  END io_product[32]
  PIN io_product[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1465.190 0.000 1465.470 4.000 ;
    END
  END io_product[33]
  PIN io_product[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1508.890 0.000 1509.170 4.000 ;
    END
  END io_product[34]
  PIN io_product[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1552.590 0.000 1552.870 4.000 ;
    END
  END io_product[35]
  PIN io_product[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1596.290 0.000 1596.570 4.000 ;
    END
  END io_product[36]
  PIN io_product[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1639.990 0.000 1640.270 4.000 ;
    END
  END io_product[37]
  PIN io_product[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1683.690 0.000 1683.970 4.000 ;
    END
  END io_product[38]
  PIN io_product[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1727.390 0.000 1727.670 4.000 ;
    END
  END io_product[39]
  PIN io_product[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END io_product[3]
  PIN io_product[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1771.090 0.000 1771.370 4.000 ;
    END
  END io_product[40]
  PIN io_product[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1814.790 0.000 1815.070 4.000 ;
    END
  END io_product[41]
  PIN io_product[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1858.490 0.000 1858.770 4.000 ;
    END
  END io_product[42]
  PIN io_product[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1902.190 0.000 1902.470 4.000 ;
    END
  END io_product[43]
  PIN io_product[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1945.890 0.000 1946.170 4.000 ;
    END
  END io_product[44]
  PIN io_product[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1989.590 0.000 1989.870 4.000 ;
    END
  END io_product[45]
  PIN io_product[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2033.290 0.000 2033.570 4.000 ;
    END
  END io_product[46]
  PIN io_product[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2076.990 0.000 2077.270 4.000 ;
    END
  END io_product[47]
  PIN io_product[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2120.690 0.000 2120.970 4.000 ;
    END
  END io_product[48]
  PIN io_product[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2164.390 0.000 2164.670 4.000 ;
    END
  END io_product[49]
  PIN io_product[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END io_product[4]
  PIN io_product[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2208.090 0.000 2208.370 4.000 ;
    END
  END io_product[50]
  PIN io_product[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2251.790 0.000 2252.070 4.000 ;
    END
  END io_product[51]
  PIN io_product[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2295.490 0.000 2295.770 4.000 ;
    END
  END io_product[52]
  PIN io_product[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2339.190 0.000 2339.470 4.000 ;
    END
  END io_product[53]
  PIN io_product[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2382.890 0.000 2383.170 4.000 ;
    END
  END io_product[54]
  PIN io_product[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2426.590 0.000 2426.870 4.000 ;
    END
  END io_product[55]
  PIN io_product[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2470.290 0.000 2470.570 4.000 ;
    END
  END io_product[56]
  PIN io_product[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2513.990 0.000 2514.270 4.000 ;
    END
  END io_product[57]
  PIN io_product[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2557.690 0.000 2557.970 4.000 ;
    END
  END io_product[58]
  PIN io_product[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2601.390 0.000 2601.670 4.000 ;
    END
  END io_product[59]
  PIN io_product[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END io_product[5]
  PIN io_product[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2645.090 0.000 2645.370 4.000 ;
    END
  END io_product[60]
  PIN io_product[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2688.790 0.000 2689.070 4.000 ;
    END
  END io_product[61]
  PIN io_product[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2732.490 0.000 2732.770 4.000 ;
    END
  END io_product[62]
  PIN io_product[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2776.190 0.000 2776.470 4.000 ;
    END
  END io_product[63]
  PIN io_product[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END io_product[6]
  PIN io_product[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END io_product[7]
  PIN io_product[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END io_product[8]
  PIN io_product[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END io_product[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.530 1756.000 2099.810 1760.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 4.670 6.840 2796.270 1749.200 ;
      LAYER met2 ;
        RECT 4.690 4.280 2796.240 1749.145 ;
        RECT 4.690 3.670 22.810 4.280 ;
        RECT 23.650 3.670 66.510 4.280 ;
        RECT 67.350 3.670 110.210 4.280 ;
        RECT 111.050 3.670 153.910 4.280 ;
        RECT 154.750 3.670 197.610 4.280 ;
        RECT 198.450 3.670 241.310 4.280 ;
        RECT 242.150 3.670 285.010 4.280 ;
        RECT 285.850 3.670 328.710 4.280 ;
        RECT 329.550 3.670 372.410 4.280 ;
        RECT 373.250 3.670 416.110 4.280 ;
        RECT 416.950 3.670 459.810 4.280 ;
        RECT 460.650 3.670 503.510 4.280 ;
        RECT 504.350 3.670 547.210 4.280 ;
        RECT 548.050 3.670 590.910 4.280 ;
        RECT 591.750 3.670 634.610 4.280 ;
        RECT 635.450 3.670 678.310 4.280 ;
        RECT 679.150 3.670 722.010 4.280 ;
        RECT 722.850 3.670 765.710 4.280 ;
        RECT 766.550 3.670 809.410 4.280 ;
        RECT 810.250 3.670 853.110 4.280 ;
        RECT 853.950 3.670 896.810 4.280 ;
        RECT 897.650 3.670 940.510 4.280 ;
        RECT 941.350 3.670 984.210 4.280 ;
        RECT 985.050 3.670 1027.910 4.280 ;
        RECT 1028.750 3.670 1071.610 4.280 ;
        RECT 1072.450 3.670 1115.310 4.280 ;
        RECT 1116.150 3.670 1159.010 4.280 ;
        RECT 1159.850 3.670 1202.710 4.280 ;
        RECT 1203.550 3.670 1246.410 4.280 ;
        RECT 1247.250 3.670 1290.110 4.280 ;
        RECT 1290.950 3.670 1333.810 4.280 ;
        RECT 1334.650 3.670 1377.510 4.280 ;
        RECT 1378.350 3.670 1421.210 4.280 ;
        RECT 1422.050 3.670 1464.910 4.280 ;
        RECT 1465.750 3.670 1508.610 4.280 ;
        RECT 1509.450 3.670 1552.310 4.280 ;
        RECT 1553.150 3.670 1596.010 4.280 ;
        RECT 1596.850 3.670 1639.710 4.280 ;
        RECT 1640.550 3.670 1683.410 4.280 ;
        RECT 1684.250 3.670 1727.110 4.280 ;
        RECT 1727.950 3.670 1770.810 4.280 ;
        RECT 1771.650 3.670 1814.510 4.280 ;
        RECT 1815.350 3.670 1858.210 4.280 ;
        RECT 1859.050 3.670 1901.910 4.280 ;
        RECT 1902.750 3.670 1945.610 4.280 ;
        RECT 1946.450 3.670 1989.310 4.280 ;
        RECT 1990.150 3.670 2033.010 4.280 ;
        RECT 2033.850 3.670 2076.710 4.280 ;
        RECT 2077.550 3.670 2120.410 4.280 ;
        RECT 2121.250 3.670 2164.110 4.280 ;
        RECT 2164.950 3.670 2207.810 4.280 ;
        RECT 2208.650 3.670 2251.510 4.280 ;
        RECT 2252.350 3.670 2295.210 4.280 ;
        RECT 2296.050 3.670 2338.910 4.280 ;
        RECT 2339.750 3.670 2382.610 4.280 ;
        RECT 2383.450 3.670 2426.310 4.280 ;
        RECT 2427.150 3.670 2470.010 4.280 ;
        RECT 2470.850 3.670 2513.710 4.280 ;
        RECT 2514.550 3.670 2557.410 4.280 ;
        RECT 2558.250 3.670 2601.110 4.280 ;
        RECT 2601.950 3.670 2644.810 4.280 ;
        RECT 2645.650 3.670 2688.510 4.280 ;
        RECT 2689.350 3.670 2732.210 4.280 ;
        RECT 2733.050 3.670 2775.910 4.280 ;
        RECT 2776.750 3.670 2796.240 4.280 ;
      LAYER met3 ;
        RECT 3.990 1722.800 2796.000 1749.125 ;
        RECT 4.400 1721.400 2795.600 1722.800 ;
        RECT 3.990 1668.400 2796.000 1721.400 ;
        RECT 4.400 1667.000 2795.600 1668.400 ;
        RECT 3.990 1614.000 2796.000 1667.000 ;
        RECT 4.400 1612.600 2795.600 1614.000 ;
        RECT 3.990 1559.600 2796.000 1612.600 ;
        RECT 4.400 1558.200 2795.600 1559.600 ;
        RECT 3.990 1505.200 2796.000 1558.200 ;
        RECT 4.400 1503.800 2795.600 1505.200 ;
        RECT 3.990 1450.800 2796.000 1503.800 ;
        RECT 4.400 1449.400 2795.600 1450.800 ;
        RECT 3.990 1396.400 2796.000 1449.400 ;
        RECT 4.400 1395.000 2795.600 1396.400 ;
        RECT 3.990 1342.000 2796.000 1395.000 ;
        RECT 4.400 1340.600 2795.600 1342.000 ;
        RECT 3.990 1287.600 2796.000 1340.600 ;
        RECT 4.400 1286.200 2795.600 1287.600 ;
        RECT 3.990 1233.200 2796.000 1286.200 ;
        RECT 4.400 1231.800 2795.600 1233.200 ;
        RECT 3.990 1178.800 2796.000 1231.800 ;
        RECT 4.400 1177.400 2795.600 1178.800 ;
        RECT 3.990 1124.400 2796.000 1177.400 ;
        RECT 4.400 1123.000 2795.600 1124.400 ;
        RECT 3.990 1070.000 2796.000 1123.000 ;
        RECT 4.400 1068.600 2795.600 1070.000 ;
        RECT 3.990 1015.600 2796.000 1068.600 ;
        RECT 4.400 1014.200 2795.600 1015.600 ;
        RECT 3.990 961.200 2796.000 1014.200 ;
        RECT 4.400 959.800 2795.600 961.200 ;
        RECT 3.990 906.800 2796.000 959.800 ;
        RECT 4.400 905.400 2795.600 906.800 ;
        RECT 3.990 852.400 2796.000 905.400 ;
        RECT 4.400 851.000 2795.600 852.400 ;
        RECT 3.990 798.000 2796.000 851.000 ;
        RECT 4.400 796.600 2795.600 798.000 ;
        RECT 3.990 743.600 2796.000 796.600 ;
        RECT 4.400 742.200 2795.600 743.600 ;
        RECT 3.990 689.200 2796.000 742.200 ;
        RECT 4.400 687.800 2795.600 689.200 ;
        RECT 3.990 634.800 2796.000 687.800 ;
        RECT 4.400 633.400 2795.600 634.800 ;
        RECT 3.990 580.400 2796.000 633.400 ;
        RECT 4.400 579.000 2795.600 580.400 ;
        RECT 3.990 526.000 2796.000 579.000 ;
        RECT 4.400 524.600 2795.600 526.000 ;
        RECT 3.990 471.600 2796.000 524.600 ;
        RECT 4.400 470.200 2795.600 471.600 ;
        RECT 3.990 417.200 2796.000 470.200 ;
        RECT 4.400 415.800 2795.600 417.200 ;
        RECT 3.990 362.800 2796.000 415.800 ;
        RECT 4.400 361.400 2795.600 362.800 ;
        RECT 3.990 308.400 2796.000 361.400 ;
        RECT 4.400 307.000 2795.600 308.400 ;
        RECT 3.990 254.000 2796.000 307.000 ;
        RECT 4.400 252.600 2795.600 254.000 ;
        RECT 3.990 199.600 2796.000 252.600 ;
        RECT 4.400 198.200 2795.600 199.600 ;
        RECT 3.990 145.200 2796.000 198.200 ;
        RECT 4.400 143.800 2795.600 145.200 ;
        RECT 3.990 90.800 2796.000 143.800 ;
        RECT 4.400 89.400 2795.600 90.800 ;
        RECT 3.990 36.400 2796.000 89.400 ;
        RECT 4.400 35.000 2795.600 36.400 ;
        RECT 3.990 8.335 2796.000 35.000 ;
      LAYER met4 ;
        RECT 1360.055 144.335 1364.985 193.625 ;
  END
END DaddaTreeMultiplier
END LIBRARY

